library verilog;
use verilog.vl_types.all;
<<<<<<< HEAD
entity \IIR_tb\ is
end \IIR_tb\;
=======
entity IIR_tb is
end IIR_tb;
>>>>>>> c6788b3
