library verilog;
use verilog.vl_types.all;
entity \IIR_tb\ is
end \IIR_tb\;
