-- -- Fiore, Neri, Ribaldone, Zheng
--
-- keyword in MAIUSCOLO (es: STD_LOGIC)
-- dati in minuscolo (es: data_in)
-- segnali di controllo in MAIUSCOLO (es: EN)
-- componenti instanziati con l'iniziale maiuscola (es: Shift_register_1)
-- i segnali attivi bassi con _n finale (es: RST_n)

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE work.all;
USE work.MBE_pkg.all;

ENTITY MBE_dadda IS
PORT(	pp_mat			: IN MATRIX_PP;
	sign_pp			: IN STD_LOGIC_VECTOR(row_pp-2 DOWNTO 0);
	data_out1		: OUT STD_LOGIC_VECTOR(2*Nb-1 DOWNTO 0);
	data_out2		: OUT STD_LOGIC_VECTOR(2*Nb-1 DOWNTO 0));
END MBE_dadda;

ARCHITECTURE structure OF MBE_dadda IS

------ COMPONENTS -------

COMPONENT FA IS 
PORT(	a,b,cin	: IN STD_LOGIC;
	s,cout	: OUT STD_LOGIC);
END COMPONENT FA;

COMPONENT HA IS 
PORT(	a,b	: IN STD_LOGIC;
	s,cout	: OUT STD_LOGIC);
END COMPONENT HA;

------ SIGNALS -------

SIGNAL mult_vmat	: VECT_MATRIX;


BEGIN


	------------------------------------------
	-- PYRAMID
	------------------------------------------

		mult_vmat(0,0)(35 DOWNTO 0) <= pp_mat(0)(35 DOWNTO 0);
		mult_vmat(0,1)(0) <= sign_pp(0);
		mult_vmat(0,1)(35 DOWNTO 2) <= pp_mat(1)(33 DOWNTO 0);
		mult_vmat(0,2)(2) <= sign_pp(1);
		mult_vmat(0,15)(36 DOWNTO 36) <= pp_mat(1)(31 DOWNTO 31);
		mult_vmat(0,2)(35 DOWNTO 4) <= pp_mat(2)(31 DOWNTO 0);
		mult_vmat(0,3)(4) <= sign_pp(2);
		mult_vmat(0,14)(38 DOWNTO 36) <= pp_mat(2)(31 DOWNTO 29);
		mult_vmat(0,3)(35 DOWNTO 6) <= pp_mat(3)(29 DOWNTO 0);
		mult_vmat(0,4)(6) <= sign_pp(3);
		mult_vmat(0,13)(40 DOWNTO 36) <= pp_mat(3)(31 DOWNTO 27);
		mult_vmat(0,4)(35 DOWNTO 8) <= pp_mat(4)(27 DOWNTO 0);
		mult_vmat(0,5)(8) <= sign_pp(4);
		mult_vmat(0,12)(42 DOWNTO 36) <= pp_mat(4)(31 DOWNTO 25);
		mult_vmat(0,5)(35 DOWNTO 10) <= pp_mat(5)(25 DOWNTO 0);
		mult_vmat(0,6)(10) <= sign_pp(5);
		mult_vmat(0,11)(44 DOWNTO 36) <= pp_mat(5)(31 DOWNTO 23);
		mult_vmat(0,6)(35 DOWNTO 12) <= pp_mat(6)(23 DOWNTO 0);
		mult_vmat(0,7)(12) <= sign_pp(6);
		mult_vmat(0,10)(46 DOWNTO 36) <= pp_mat(6)(31 DOWNTO 21);
		mult_vmat(0,7)(35 DOWNTO 14) <= pp_mat(7)(21 DOWNTO 0);
		mult_vmat(0,8)(14) <= sign_pp(7);
		mult_vmat(0,9)(48 DOWNTO 36) <= pp_mat(7)(31 DOWNTO 19);
		mult_vmat(0,8)(35 DOWNTO 16) <= pp_mat(8)(19 DOWNTO 0);
		mult_vmat(0,9)(16) <= sign_pp(8);
		mult_vmat(0,8)(50 DOWNTO 36) <= pp_mat(8)(31 DOWNTO 17);
		mult_vmat(0,9)(35 DOWNTO 18) <= pp_mat(9)(17 DOWNTO 0);
		mult_vmat(0,10)(18) <= sign_pp(9);
		mult_vmat(0,7)(52 DOWNTO 36) <= pp_mat(9)(31 DOWNTO 15);
		mult_vmat(0,10)(35 DOWNTO 20) <= pp_mat(10)(15 DOWNTO 0);
		mult_vmat(0,11)(20) <= sign_pp(10);
		mult_vmat(0,6)(54 DOWNTO 36) <= pp_mat(10)(31 DOWNTO 13);
		mult_vmat(0,11)(35 DOWNTO 22) <= pp_mat(11)(13 DOWNTO 0);
		mult_vmat(0,12)(22) <= sign_pp(11);
		mult_vmat(0,5)(56 DOWNTO 36) <= pp_mat(11)(31 DOWNTO 11);
		mult_vmat(0,12)(35 DOWNTO 24) <= pp_mat(12)(11 DOWNTO 0);
		mult_vmat(0,13)(24) <= sign_pp(12);
		mult_vmat(0,4)(58 DOWNTO 36) <= pp_mat(12)(31 DOWNTO 9);
		mult_vmat(0,13)(35 DOWNTO 26) <= pp_mat(13)(9 DOWNTO 0);
		mult_vmat(0,14)(26) <= sign_pp(13);
		mult_vmat(0,3)(60 DOWNTO 36) <= pp_mat(13)(31 DOWNTO 7);
		mult_vmat(0,14)(35 DOWNTO 28) <= pp_mat(14)(7 DOWNTO 0);
		mult_vmat(0,15)(28) <= sign_pp(14);
		mult_vmat(0,2)(62 DOWNTO 36) <= pp_mat(14)(31 DOWNTO 5);
		mult_vmat(0,15)(35 DOWNTO 30) <= pp_mat(15)(5 DOWNTO 0);
		mult_vmat(0,16)(30) <= sign_pp(15);
		mult_vmat(0,1)(63 DOWNTO 36) <= pp_mat(15)(30 DOWNTO 3);
		mult_vmat(0,16)(35 DOWNTO 32) <= pp_mat(16)(3 DOWNTO 0);
		mult_vmat(0,0)(63 DOWNTO 36) <= pp_mat(16)(28 DOWNTO 1);


	------------------------------------------
	-- LEVEL 1
	------------------------------------------


		-- COLUMN 1
		mult_vmat(1,0)(0) <= mult_vmat(0,0)(0);
		mult_vmat(1,1)(0) <= mult_vmat(0,1)(0);

		-- COLUMN 2
		mult_vmat(1,0)(1) <= mult_vmat(0,0)(1);

		-- COLUMN 3
		mult_vmat(1,0)(2) <= mult_vmat(0,0)(2);
		mult_vmat(1,1)(2) <= mult_vmat(0,1)(2);
		mult_vmat(1,2)(2) <= mult_vmat(0,2)(2);

		-- COLUMN 4
		mult_vmat(1,0)(3) <= mult_vmat(0,0)(3);
		mult_vmat(1,1)(3) <= mult_vmat(0,1)(3);

		-- COLUMN 5
		mult_vmat(1,0)(4) <= mult_vmat(0,0)(4);
		mult_vmat(1,1)(4) <= mult_vmat(0,1)(4);
		mult_vmat(1,2)(4) <= mult_vmat(0,2)(4);
		mult_vmat(1,3)(4) <= mult_vmat(0,3)(4);

		-- COLUMN 6
		mult_vmat(1,0)(5) <= mult_vmat(0,0)(5);
		mult_vmat(1,1)(5) <= mult_vmat(0,1)(5);
		mult_vmat(1,2)(5) <= mult_vmat(0,2)(5);

		-- COLUMN 7
		mult_vmat(1,0)(6) <= mult_vmat(0,0)(6);
		mult_vmat(1,1)(6) <= mult_vmat(0,1)(6);
		mult_vmat(1,2)(6) <= mult_vmat(0,2)(6);
		mult_vmat(1,3)(6) <= mult_vmat(0,3)(6);
		mult_vmat(1,4)(6) <= mult_vmat(0,4)(6);

		-- COLUMN 8
		mult_vmat(1,0)(7) <= mult_vmat(0,0)(7);
		mult_vmat(1,1)(7) <= mult_vmat(0,1)(7);
		mult_vmat(1,2)(7) <= mult_vmat(0,2)(7);
		mult_vmat(1,3)(7) <= mult_vmat(0,3)(7);

		-- COLUMN 9
		mult_vmat(1,0)(8) <= mult_vmat(0,0)(8);
		mult_vmat(1,1)(8) <= mult_vmat(0,1)(8);
		mult_vmat(1,2)(8) <= mult_vmat(0,2)(8);
		mult_vmat(1,3)(8) <= mult_vmat(0,3)(8);
		mult_vmat(1,4)(8) <= mult_vmat(0,4)(8);
		mult_vmat(1,5)(8) <= mult_vmat(0,5)(8);

		-- COLUMN 10
		mult_vmat(1,0)(9) <= mult_vmat(0,0)(9);
		mult_vmat(1,1)(9) <= mult_vmat(0,1)(9);
		mult_vmat(1,2)(9) <= mult_vmat(0,2)(9);
		mult_vmat(1,3)(9) <= mult_vmat(0,3)(9);
		mult_vmat(1,4)(9) <= mult_vmat(0,4)(9);

		-- COLUMN 11
		mult_vmat(1,0)(10) <= mult_vmat(0,0)(10);
		mult_vmat(1,1)(10) <= mult_vmat(0,1)(10);
		mult_vmat(1,2)(10) <= mult_vmat(0,2)(10);
		mult_vmat(1,3)(10) <= mult_vmat(0,3)(10);
		mult_vmat(1,4)(10) <= mult_vmat(0,4)(10);
		mult_vmat(1,5)(10) <= mult_vmat(0,5)(10);
		mult_vmat(1,6)(10) <= mult_vmat(0,6)(10);

		-- COLUMN 12
		mult_vmat(1,0)(11) <= mult_vmat(0,0)(11);
		mult_vmat(1,1)(11) <= mult_vmat(0,1)(11);
		mult_vmat(1,2)(11) <= mult_vmat(0,2)(11);
		mult_vmat(1,3)(11) <= mult_vmat(0,3)(11);
		mult_vmat(1,4)(11) <= mult_vmat(0,4)(11);
		mult_vmat(1,5)(11) <= mult_vmat(0,5)(11);

		-- COLUMN 13
		mult_vmat(1,0)(12) <= mult_vmat(0,0)(12);
		mult_vmat(1,1)(12) <= mult_vmat(0,1)(12);
		mult_vmat(1,2)(12) <= mult_vmat(0,2)(12);
		mult_vmat(1,3)(12) <= mult_vmat(0,3)(12);
		mult_vmat(1,4)(12) <= mult_vmat(0,4)(12);
		mult_vmat(1,5)(12) <= mult_vmat(0,5)(12);
		mult_vmat(1,6)(12) <= mult_vmat(0,6)(12);
		mult_vmat(1,7)(12) <= mult_vmat(0,7)(12);

		-- COLUMN 14
		mult_vmat(1,0)(13) <= mult_vmat(0,0)(13);
		mult_vmat(1,1)(13) <= mult_vmat(0,1)(13);
		mult_vmat(1,2)(13) <= mult_vmat(0,2)(13);
		mult_vmat(1,3)(13) <= mult_vmat(0,3)(13);
		mult_vmat(1,4)(13) <= mult_vmat(0,4)(13);
		mult_vmat(1,5)(13) <= mult_vmat(0,5)(13);
		mult_vmat(1,6)(13) <= mult_vmat(0,6)(13);

		-- COLUMN 15
		mult_vmat(1,0)(14) <= mult_vmat(0,0)(14);
		mult_vmat(1,1)(14) <= mult_vmat(0,1)(14);
		mult_vmat(1,2)(14) <= mult_vmat(0,2)(14);
		mult_vmat(1,3)(14) <= mult_vmat(0,3)(14);
		mult_vmat(1,4)(14) <= mult_vmat(0,4)(14);
		mult_vmat(1,5)(14) <= mult_vmat(0,5)(14);
		mult_vmat(1,6)(14) <= mult_vmat(0,6)(14);
		mult_vmat(1,7)(14) <= mult_vmat(0,7)(14);
		mult_vmat(1,8)(14) <= mult_vmat(0,8)(14);

		-- COLUMN 16
		mult_vmat(1,0)(15) <= mult_vmat(0,0)(15);
		mult_vmat(1,1)(15) <= mult_vmat(0,1)(15);
		mult_vmat(1,2)(15) <= mult_vmat(0,2)(15);
		mult_vmat(1,3)(15) <= mult_vmat(0,3)(15);
		mult_vmat(1,4)(15) <= mult_vmat(0,4)(15);
		mult_vmat(1,5)(15) <= mult_vmat(0,5)(15);
		mult_vmat(1,6)(15) <= mult_vmat(0,6)(15);
		mult_vmat(1,7)(15) <= mult_vmat(0,7)(15);

		-- COLUMN 17
		mult_vmat(1,0)(16) <= mult_vmat(0,0)(16);
		mult_vmat(1,1)(16) <= mult_vmat(0,1)(16);
		mult_vmat(1,2)(16) <= mult_vmat(0,2)(16);
		mult_vmat(1,3)(16) <= mult_vmat(0,3)(16);
		mult_vmat(1,4)(16) <= mult_vmat(0,4)(16);
		mult_vmat(1,5)(16) <= mult_vmat(0,5)(16);
		mult_vmat(1,6)(16) <= mult_vmat(0,6)(16);
		mult_vmat(1,7)(16) <= mult_vmat(0,7)(16);
		mult_vmat(1,8)(16) <= mult_vmat(0,8)(16);
		mult_vmat(1,9)(16) <= mult_vmat(0,9)(16);

		-- COLUMN 18
		mult_vmat(1,0)(17) <= mult_vmat(0,0)(17);
		mult_vmat(1,1)(17) <= mult_vmat(0,1)(17);
		mult_vmat(1,2)(17) <= mult_vmat(0,2)(17);
		mult_vmat(1,3)(17) <= mult_vmat(0,3)(17);
		mult_vmat(1,4)(17) <= mult_vmat(0,4)(17);
		mult_vmat(1,5)(17) <= mult_vmat(0,5)(17);
		mult_vmat(1,6)(17) <= mult_vmat(0,6)(17);
		mult_vmat(1,7)(17) <= mult_vmat(0,7)(17);
		mult_vmat(1,8)(17) <= mult_vmat(0,8)(17);

		-- COLUMN 19
		mult_vmat(1,0)(18) <= mult_vmat(0,0)(18);
		mult_vmat(1,1)(18) <= mult_vmat(0,1)(18);
		mult_vmat(1,2)(18) <= mult_vmat(0,2)(18);
		mult_vmat(1,3)(18) <= mult_vmat(0,3)(18);
		mult_vmat(1,4)(18) <= mult_vmat(0,4)(18);
		mult_vmat(1,5)(18) <= mult_vmat(0,5)(18);
		mult_vmat(1,6)(18) <= mult_vmat(0,6)(18);
		mult_vmat(1,7)(18) <= mult_vmat(0,7)(18);
		mult_vmat(1,8)(18) <= mult_vmat(0,8)(18);
		mult_vmat(1,9)(18) <= mult_vmat(0,9)(18);
		mult_vmat(1,10)(18) <= mult_vmat(0,10)(18);

		-- COLUMN 20
		mult_vmat(1,0)(19) <= mult_vmat(0,0)(19);
		mult_vmat(1,1)(19) <= mult_vmat(0,1)(19);
		mult_vmat(1,2)(19) <= mult_vmat(0,2)(19);
		mult_vmat(1,3)(19) <= mult_vmat(0,3)(19);
		mult_vmat(1,4)(19) <= mult_vmat(0,4)(19);
		mult_vmat(1,5)(19) <= mult_vmat(0,5)(19);
		mult_vmat(1,6)(19) <= mult_vmat(0,6)(19);
		mult_vmat(1,7)(19) <= mult_vmat(0,7)(19);
		mult_vmat(1,8)(19) <= mult_vmat(0,8)(19);
		mult_vmat(1,9)(19) <= mult_vmat(0,9)(19);

		-- COLUMN 21
		mult_vmat(1,0)(20) <= mult_vmat(0,0)(20);
		mult_vmat(1,1)(20) <= mult_vmat(0,1)(20);
		mult_vmat(1,2)(20) <= mult_vmat(0,2)(20);
		mult_vmat(1,3)(20) <= mult_vmat(0,3)(20);
		mult_vmat(1,4)(20) <= mult_vmat(0,4)(20);
		mult_vmat(1,5)(20) <= mult_vmat(0,5)(20);
		mult_vmat(1,6)(20) <= mult_vmat(0,6)(20);
		mult_vmat(1,7)(20) <= mult_vmat(0,7)(20);
		mult_vmat(1,8)(20) <= mult_vmat(0,8)(20);
		mult_vmat(1,9)(20) <= mult_vmat(0,9)(20);
		mult_vmat(1,10)(20) <= mult_vmat(0,10)(20);
		mult_vmat(1,11)(20) <= mult_vmat(0,11)(20);

		-- COLUMN 22
		mult_vmat(1,0)(21) <= mult_vmat(0,0)(21);
		mult_vmat(1,1)(21) <= mult_vmat(0,1)(21);
		mult_vmat(1,2)(21) <= mult_vmat(0,2)(21);
		mult_vmat(1,3)(21) <= mult_vmat(0,3)(21);
		mult_vmat(1,4)(21) <= mult_vmat(0,4)(21);
		mult_vmat(1,5)(21) <= mult_vmat(0,5)(21);
		mult_vmat(1,6)(21) <= mult_vmat(0,6)(21);
		mult_vmat(1,7)(21) <= mult_vmat(0,7)(21);
		mult_vmat(1,8)(21) <= mult_vmat(0,8)(21);
		mult_vmat(1,9)(21) <= mult_vmat(0,9)(21);
		mult_vmat(1,10)(21) <= mult_vmat(0,10)(21);

		-- COLUMN 23
		mult_vmat(1,0)(22) <= mult_vmat(0,0)(22);
		mult_vmat(1,1)(22) <= mult_vmat(0,1)(22);
		mult_vmat(1,2)(22) <= mult_vmat(0,2)(22);
		mult_vmat(1,3)(22) <= mult_vmat(0,3)(22);
		mult_vmat(1,4)(22) <= mult_vmat(0,4)(22);
		mult_vmat(1,5)(22) <= mult_vmat(0,5)(22);
		mult_vmat(1,6)(22) <= mult_vmat(0,6)(22);
		mult_vmat(1,7)(22) <= mult_vmat(0,7)(22);
		mult_vmat(1,8)(22) <= mult_vmat(0,8)(22);
		mult_vmat(1,9)(22) <= mult_vmat(0,9)(22);
		mult_vmat(1,10)(22) <= mult_vmat(0,10)(22);
		mult_vmat(1,11)(22) <= mult_vmat(0,11)(22);
		mult_vmat(1,12)(22) <= mult_vmat(0,12)(22);

		-- COLUMN 24
		mult_vmat(1,0)(23) <= mult_vmat(0,0)(23);
		mult_vmat(1,1)(23) <= mult_vmat(0,1)(23);
		mult_vmat(1,2)(23) <= mult_vmat(0,2)(23);
		mult_vmat(1,3)(23) <= mult_vmat(0,3)(23);
		mult_vmat(1,4)(23) <= mult_vmat(0,4)(23);
		mult_vmat(1,5)(23) <= mult_vmat(0,5)(23);
		mult_vmat(1,6)(23) <= mult_vmat(0,6)(23);
		mult_vmat(1,7)(23) <= mult_vmat(0,7)(23);
		mult_vmat(1,8)(23) <= mult_vmat(0,8)(23);
		mult_vmat(1,9)(23) <= mult_vmat(0,9)(23);
		mult_vmat(1,10)(23) <= mult_vmat(0,10)(23);
		mult_vmat(1,11)(23) <= mult_vmat(0,11)(23);

		-- COLUMN 25

		HA_0_24: HA PORT MAP (
			mult_vmat(0,0)(24),
			mult_vmat(0,1)(24),
			mult_vmat(1,0)(24),
			mult_vmat(1,0)(25)
		);

		mult_vmat(1,1)(24) <= mult_vmat(0,2)(24);
		mult_vmat(1,2)(24) <= mult_vmat(0,3)(24);
		mult_vmat(1,3)(24) <= mult_vmat(0,4)(24);
		mult_vmat(1,4)(24) <= mult_vmat(0,5)(24);
		mult_vmat(1,5)(24) <= mult_vmat(0,6)(24);
		mult_vmat(1,6)(24) <= mult_vmat(0,7)(24);
		mult_vmat(1,7)(24) <= mult_vmat(0,8)(24);
		mult_vmat(1,8)(24) <= mult_vmat(0,9)(24);
		mult_vmat(1,9)(24) <= mult_vmat(0,10)(24);
		mult_vmat(1,10)(24) <= mult_vmat(0,11)(24);
		mult_vmat(1,11)(24) <= mult_vmat(0,12)(24);
		mult_vmat(1,12)(24) <= mult_vmat(0,13)(24);

		-- COLUMN 26

		HA_0_25: HA PORT MAP (
			mult_vmat(0,0)(25),
			mult_vmat(0,1)(25),
			mult_vmat(1,1)(25),
			mult_vmat(1,0)(26)
		);

		mult_vmat(1,2)(25) <= mult_vmat(0,2)(25);
		mult_vmat(1,3)(25) <= mult_vmat(0,3)(25);
		mult_vmat(1,4)(25) <= mult_vmat(0,4)(25);
		mult_vmat(1,5)(25) <= mult_vmat(0,5)(25);
		mult_vmat(1,6)(25) <= mult_vmat(0,6)(25);
		mult_vmat(1,7)(25) <= mult_vmat(0,7)(25);
		mult_vmat(1,8)(25) <= mult_vmat(0,8)(25);
		mult_vmat(1,9)(25) <= mult_vmat(0,9)(25);
		mult_vmat(1,10)(25) <= mult_vmat(0,10)(25);
		mult_vmat(1,11)(25) <= mult_vmat(0,11)(25);
		mult_vmat(1,12)(25) <= mult_vmat(0,12)(25);

		-- COLUMN 27

		FA_0_26_1: FA PORT MAP (
			mult_vmat(0,0)(26),
			mult_vmat(0,1)(26),
			mult_vmat(0,2)(26),
			mult_vmat(1,1)(26),
			mult_vmat(1,0)(27)
		);


		HA_0_26: HA PORT MAP (
			mult_vmat(0,3)(26),
			mult_vmat(0,4)(26),
			mult_vmat(1,2)(26),
			mult_vmat(1,1)(27)
		);

		mult_vmat(1,3)(26) <= mult_vmat(0,5)(26);
		mult_vmat(1,4)(26) <= mult_vmat(0,6)(26);
		mult_vmat(1,5)(26) <= mult_vmat(0,7)(26);
		mult_vmat(1,6)(26) <= mult_vmat(0,8)(26);
		mult_vmat(1,7)(26) <= mult_vmat(0,9)(26);
		mult_vmat(1,8)(26) <= mult_vmat(0,10)(26);
		mult_vmat(1,9)(26) <= mult_vmat(0,11)(26);
		mult_vmat(1,10)(26) <= mult_vmat(0,12)(26);
		mult_vmat(1,11)(26) <= mult_vmat(0,13)(26);
		mult_vmat(1,12)(26) <= mult_vmat(0,14)(26);

		-- COLUMN 28

		FA_0_27_1: FA PORT MAP (
			mult_vmat(0,0)(27),
			mult_vmat(0,1)(27),
			mult_vmat(0,2)(27),
			mult_vmat(1,2)(27),
			mult_vmat(1,0)(28)
		);


		HA_0_27: HA PORT MAP (
			mult_vmat(0,3)(27),
			mult_vmat(0,4)(27),
			mult_vmat(1,3)(27),
			mult_vmat(1,1)(28)
		);

		mult_vmat(1,4)(27) <= mult_vmat(0,5)(27);
		mult_vmat(1,5)(27) <= mult_vmat(0,6)(27);
		mult_vmat(1,6)(27) <= mult_vmat(0,7)(27);
		mult_vmat(1,7)(27) <= mult_vmat(0,8)(27);
		mult_vmat(1,8)(27) <= mult_vmat(0,9)(27);
		mult_vmat(1,9)(27) <= mult_vmat(0,10)(27);
		mult_vmat(1,10)(27) <= mult_vmat(0,11)(27);
		mult_vmat(1,11)(27) <= mult_vmat(0,12)(27);
		mult_vmat(1,12)(27) <= mult_vmat(0,13)(27);

		-- COLUMN 29

		FA_0_28_1: FA PORT MAP (
			mult_vmat(0,0)(28),
			mult_vmat(0,1)(28),
			mult_vmat(0,2)(28),
			mult_vmat(1,2)(28),
			mult_vmat(1,0)(29)
		);


		FA_0_28_2: FA PORT MAP (
			mult_vmat(0,3)(28),
			mult_vmat(0,4)(28),
			mult_vmat(0,5)(28),
			mult_vmat(1,3)(28),
			mult_vmat(1,1)(29)
		);


		HA_0_28: HA PORT MAP (
			mult_vmat(0,6)(28),
			mult_vmat(0,7)(28),
			mult_vmat(1,4)(28),
			mult_vmat(1,2)(29)
		);

		mult_vmat(1,5)(28) <= mult_vmat(0,8)(28);
		mult_vmat(1,6)(28) <= mult_vmat(0,9)(28);
		mult_vmat(1,7)(28) <= mult_vmat(0,10)(28);
		mult_vmat(1,8)(28) <= mult_vmat(0,11)(28);
		mult_vmat(1,9)(28) <= mult_vmat(0,12)(28);
		mult_vmat(1,10)(28) <= mult_vmat(0,13)(28);
		mult_vmat(1,11)(28) <= mult_vmat(0,14)(28);
		mult_vmat(1,12)(28) <= mult_vmat(0,15)(28);

		-- COLUMN 30

		FA_0_29_1: FA PORT MAP (
			mult_vmat(0,0)(29),
			mult_vmat(0,1)(29),
			mult_vmat(0,2)(29),
			mult_vmat(1,3)(29),
			mult_vmat(1,0)(30)
		);


		FA_0_29_2: FA PORT MAP (
			mult_vmat(0,3)(29),
			mult_vmat(0,4)(29),
			mult_vmat(0,5)(29),
			mult_vmat(1,4)(29),
			mult_vmat(1,1)(30)
		);


		HA_0_29: HA PORT MAP (
			mult_vmat(0,6)(29),
			mult_vmat(0,7)(29),
			mult_vmat(1,5)(29),
			mult_vmat(1,2)(30)
		);

		mult_vmat(1,6)(29) <= mult_vmat(0,8)(29);
		mult_vmat(1,7)(29) <= mult_vmat(0,9)(29);
		mult_vmat(1,8)(29) <= mult_vmat(0,10)(29);
		mult_vmat(1,9)(29) <= mult_vmat(0,11)(29);
		mult_vmat(1,10)(29) <= mult_vmat(0,12)(29);
		mult_vmat(1,11)(29) <= mult_vmat(0,13)(29);
		mult_vmat(1,12)(29) <= mult_vmat(0,14)(29);

		-- COLUMN 31

		FA_0_30_1: FA PORT MAP (
			mult_vmat(0,0)(30),
			mult_vmat(0,1)(30),
			mult_vmat(0,2)(30),
			mult_vmat(1,3)(30),
			mult_vmat(1,0)(31)
		);


		FA_0_30_2: FA PORT MAP (
			mult_vmat(0,3)(30),
			mult_vmat(0,4)(30),
			mult_vmat(0,5)(30),
			mult_vmat(1,4)(30),
			mult_vmat(1,1)(31)
		);


		FA_0_30_3: FA PORT MAP (
			mult_vmat(0,6)(30),
			mult_vmat(0,7)(30),
			mult_vmat(0,8)(30),
			mult_vmat(1,5)(30),
			mult_vmat(1,2)(31)
		);


		HA_0_30: HA PORT MAP (
			mult_vmat(0,9)(30),
			mult_vmat(0,10)(30),
			mult_vmat(1,6)(30),
			mult_vmat(1,3)(31)
		);

		mult_vmat(1,7)(30) <= mult_vmat(0,11)(30);
		mult_vmat(1,8)(30) <= mult_vmat(0,12)(30);
		mult_vmat(1,9)(30) <= mult_vmat(0,13)(30);
		mult_vmat(1,10)(30) <= mult_vmat(0,14)(30);
		mult_vmat(1,11)(30) <= mult_vmat(0,15)(30);
		mult_vmat(1,12)(30) <= mult_vmat(0,16)(30);

		-- COLUMN 32

		FA_0_31_1: FA PORT MAP (
			mult_vmat(0,0)(31),
			mult_vmat(0,1)(31),
			mult_vmat(0,2)(31),
			mult_vmat(1,4)(31),
			mult_vmat(1,0)(32)
		);


		FA_0_31_2: FA PORT MAP (
			mult_vmat(0,3)(31),
			mult_vmat(0,4)(31),
			mult_vmat(0,5)(31),
			mult_vmat(1,5)(31),
			mult_vmat(1,1)(32)
		);


		FA_0_31_3: FA PORT MAP (
			mult_vmat(0,6)(31),
			mult_vmat(0,7)(31),
			mult_vmat(0,8)(31),
			mult_vmat(1,6)(31),
			mult_vmat(1,2)(32)
		);


		HA_0_31: HA PORT MAP (
			mult_vmat(0,9)(31),
			mult_vmat(0,10)(31),
			mult_vmat(1,7)(31),
			mult_vmat(1,3)(32)
		);

		mult_vmat(1,8)(31) <= mult_vmat(0,11)(31);
		mult_vmat(1,9)(31) <= mult_vmat(0,12)(31);
		mult_vmat(1,10)(31) <= mult_vmat(0,13)(31);
		mult_vmat(1,11)(31) <= mult_vmat(0,14)(31);
		mult_vmat(1,12)(31) <= mult_vmat(0,15)(31);

		-- COLUMN 33

		FA_0_32_1: FA PORT MAP (
			mult_vmat(0,0)(32),
			mult_vmat(0,1)(32),
			mult_vmat(0,2)(32),
			mult_vmat(1,4)(32),
			mult_vmat(1,0)(33)
		);


		FA_0_32_2: FA PORT MAP (
			mult_vmat(0,3)(32),
			mult_vmat(0,4)(32),
			mult_vmat(0,5)(32),
			mult_vmat(1,5)(32),
			mult_vmat(1,1)(33)
		);


		FA_0_32_3: FA PORT MAP (
			mult_vmat(0,6)(32),
			mult_vmat(0,7)(32),
			mult_vmat(0,8)(32),
			mult_vmat(1,6)(32),
			mult_vmat(1,2)(33)
		);


		FA_0_32_4: FA PORT MAP (
			mult_vmat(0,9)(32),
			mult_vmat(0,10)(32),
			mult_vmat(0,11)(32),
			mult_vmat(1,7)(32),
			mult_vmat(1,3)(33)
		);

		mult_vmat(1,8)(32) <= mult_vmat(0,12)(32);
		mult_vmat(1,9)(32) <= mult_vmat(0,13)(32);
		mult_vmat(1,10)(32) <= mult_vmat(0,14)(32);
		mult_vmat(1,11)(32) <= mult_vmat(0,15)(32);
		mult_vmat(1,12)(32) <= mult_vmat(0,16)(32);

		-- COLUMN 34

		FA_0_33_1: FA PORT MAP (
			mult_vmat(0,0)(33),
			mult_vmat(0,1)(33),
			mult_vmat(0,2)(33),
			mult_vmat(1,4)(33),
			mult_vmat(1,0)(34)
		);


		FA_0_33_2: FA PORT MAP (
			mult_vmat(0,3)(33),
			mult_vmat(0,4)(33),
			mult_vmat(0,5)(33),
			mult_vmat(1,5)(33),
			mult_vmat(1,1)(34)
		);


		FA_0_33_3: FA PORT MAP (
			mult_vmat(0,6)(33),
			mult_vmat(0,7)(33),
			mult_vmat(0,8)(33),
			mult_vmat(1,6)(33),
			mult_vmat(1,2)(34)
		);


		FA_0_33_4: FA PORT MAP (
			mult_vmat(0,9)(33),
			mult_vmat(0,10)(33),
			mult_vmat(0,11)(33),
			mult_vmat(1,7)(33),
			mult_vmat(1,3)(34)
		);

		mult_vmat(1,8)(33) <= mult_vmat(0,12)(33);
		mult_vmat(1,9)(33) <= mult_vmat(0,13)(33);
		mult_vmat(1,10)(33) <= mult_vmat(0,14)(33);
		mult_vmat(1,11)(33) <= mult_vmat(0,15)(33);
		mult_vmat(1,12)(33) <= mult_vmat(0,16)(33);

		-- COLUMN 35

		FA_0_34_1: FA PORT MAP (
			mult_vmat(0,0)(34),
			mult_vmat(0,1)(34),
			mult_vmat(0,2)(34),
			mult_vmat(1,4)(34),
			mult_vmat(1,0)(35)
		);


		FA_0_34_2: FA PORT MAP (
			mult_vmat(0,3)(34),
			mult_vmat(0,4)(34),
			mult_vmat(0,5)(34),
			mult_vmat(1,5)(34),
			mult_vmat(1,1)(35)
		);


		FA_0_34_3: FA PORT MAP (
			mult_vmat(0,6)(34),
			mult_vmat(0,7)(34),
			mult_vmat(0,8)(34),
			mult_vmat(1,6)(34),
			mult_vmat(1,2)(35)
		);


		FA_0_34_4: FA PORT MAP (
			mult_vmat(0,9)(34),
			mult_vmat(0,10)(34),
			mult_vmat(0,11)(34),
			mult_vmat(1,7)(34),
			mult_vmat(1,3)(35)
		);

		mult_vmat(1,8)(34) <= mult_vmat(0,12)(34);
		mult_vmat(1,9)(34) <= mult_vmat(0,13)(34);
		mult_vmat(1,10)(34) <= mult_vmat(0,14)(34);
		mult_vmat(1,11)(34) <= mult_vmat(0,15)(34);
		mult_vmat(1,12)(34) <= mult_vmat(0,16)(34);

		-- COLUMN 36

		FA_0_35_1: FA PORT MAP (
			mult_vmat(0,0)(35),
			mult_vmat(0,1)(35),
			mult_vmat(0,2)(35),
			mult_vmat(1,4)(35),
			mult_vmat(1,0)(36)
		);


		FA_0_35_2: FA PORT MAP (
			mult_vmat(0,3)(35),
			mult_vmat(0,4)(35),
			mult_vmat(0,5)(35),
			mult_vmat(1,5)(35),
			mult_vmat(1,1)(36)
		);


		FA_0_35_3: FA PORT MAP (
			mult_vmat(0,6)(35),
			mult_vmat(0,7)(35),
			mult_vmat(0,8)(35),
			mult_vmat(1,6)(35),
			mult_vmat(1,2)(36)
		);


		FA_0_35_4: FA PORT MAP (
			mult_vmat(0,9)(35),
			mult_vmat(0,10)(35),
			mult_vmat(0,11)(35),
			mult_vmat(1,7)(35),
			mult_vmat(1,3)(36)
		);

		mult_vmat(1,8)(35) <= mult_vmat(0,12)(35);
		mult_vmat(1,9)(35) <= mult_vmat(0,13)(35);
		mult_vmat(1,10)(35) <= mult_vmat(0,14)(35);
		mult_vmat(1,11)(35) <= mult_vmat(0,15)(35);
		mult_vmat(1,12)(35) <= mult_vmat(0,16)(35);

		-- COLUMN 37

		FA_0_36_1: FA PORT MAP (
			mult_vmat(0,0)(36),
			mult_vmat(0,1)(36),
			mult_vmat(0,2)(36),
			mult_vmat(1,4)(36),
			mult_vmat(1,0)(37)
		);


		FA_0_36_2: FA PORT MAP (
			mult_vmat(0,3)(36),
			mult_vmat(0,4)(36),
			mult_vmat(0,5)(36),
			mult_vmat(1,5)(36),
			mult_vmat(1,1)(37)
		);


		FA_0_36_3: FA PORT MAP (
			mult_vmat(0,6)(36),
			mult_vmat(0,7)(36),
			mult_vmat(0,8)(36),
			mult_vmat(1,6)(36),
			mult_vmat(1,2)(37)
		);


		HA_0_36: HA PORT MAP (
			mult_vmat(0,9)(36),
			mult_vmat(0,10)(36),
			mult_vmat(1,7)(36),
			mult_vmat(1,3)(37)
		);

		mult_vmat(1,8)(36) <= mult_vmat(0,11)(36);
		mult_vmat(1,9)(36) <= mult_vmat(0,12)(36);
		mult_vmat(1,10)(36) <= mult_vmat(0,13)(36);
		mult_vmat(1,11)(36) <= mult_vmat(0,14)(36);
		mult_vmat(1,12)(36) <= mult_vmat(0,15)(36);

		-- COLUMN 38

		FA_0_37_1: FA PORT MAP (
			mult_vmat(0,0)(37),
			mult_vmat(0,1)(37),
			mult_vmat(0,2)(37),
			mult_vmat(1,4)(37),
			mult_vmat(1,0)(38)
		);


		FA_0_37_2: FA PORT MAP (
			mult_vmat(0,3)(37),
			mult_vmat(0,4)(37),
			mult_vmat(0,5)(37),
			mult_vmat(1,5)(37),
			mult_vmat(1,1)(38)
		);


		FA_0_37_3: FA PORT MAP (
			mult_vmat(0,6)(37),
			mult_vmat(0,7)(37),
			mult_vmat(0,8)(37),
			mult_vmat(1,6)(37),
			mult_vmat(1,2)(38)
		);

		mult_vmat(1,7)(37) <= mult_vmat(0,9)(37);
		mult_vmat(1,8)(37) <= mult_vmat(0,10)(37);
		mult_vmat(1,9)(37) <= mult_vmat(0,11)(37);
		mult_vmat(1,10)(37) <= mult_vmat(0,12)(37);
		mult_vmat(1,11)(37) <= mult_vmat(0,13)(37);
		mult_vmat(1,12)(37) <= mult_vmat(0,14)(37);

		-- COLUMN 39

		FA_0_38_1: FA PORT MAP (
			mult_vmat(0,0)(38),
			mult_vmat(0,1)(38),
			mult_vmat(0,2)(38),
			mult_vmat(1,3)(38),
			mult_vmat(1,0)(39)
		);


		FA_0_38_2: FA PORT MAP (
			mult_vmat(0,3)(38),
			mult_vmat(0,4)(38),
			mult_vmat(0,5)(38),
			mult_vmat(1,4)(38),
			mult_vmat(1,1)(39)
		);


		HA_0_38: HA PORT MAP (
			mult_vmat(0,6)(38),
			mult_vmat(0,7)(38),
			mult_vmat(1,5)(38),
			mult_vmat(1,2)(39)
		);

		mult_vmat(1,6)(38) <= mult_vmat(0,8)(38);
		mult_vmat(1,7)(38) <= mult_vmat(0,9)(38);
		mult_vmat(1,8)(38) <= mult_vmat(0,10)(38);
		mult_vmat(1,9)(38) <= mult_vmat(0,11)(38);
		mult_vmat(1,10)(38) <= mult_vmat(0,12)(38);
		mult_vmat(1,11)(38) <= mult_vmat(0,13)(38);
		mult_vmat(1,12)(38) <= mult_vmat(0,14)(38);

		-- COLUMN 40

		FA_0_39_1: FA PORT MAP (
			mult_vmat(0,0)(39),
			mult_vmat(0,1)(39),
			mult_vmat(0,2)(39),
			mult_vmat(1,3)(39),
			mult_vmat(1,0)(40)
		);


		FA_0_39_2: FA PORT MAP (
			mult_vmat(0,3)(39),
			mult_vmat(0,4)(39),
			mult_vmat(0,5)(39),
			mult_vmat(1,4)(39),
			mult_vmat(1,1)(40)
		);

		mult_vmat(1,5)(39) <= mult_vmat(0,6)(39);
		mult_vmat(1,6)(39) <= mult_vmat(0,7)(39);
		mult_vmat(1,7)(39) <= mult_vmat(0,8)(39);
		mult_vmat(1,8)(39) <= mult_vmat(0,9)(39);
		mult_vmat(1,9)(39) <= mult_vmat(0,10)(39);
		mult_vmat(1,10)(39) <= mult_vmat(0,11)(39);
		mult_vmat(1,11)(39) <= mult_vmat(0,12)(39);
		mult_vmat(1,12)(39) <= mult_vmat(0,13)(39);

		-- COLUMN 41

		FA_0_40_1: FA PORT MAP (
			mult_vmat(0,0)(40),
			mult_vmat(0,1)(40),
			mult_vmat(0,2)(40),
			mult_vmat(1,2)(40),
			mult_vmat(1,0)(41)
		);


		HA_0_40: HA PORT MAP (
			mult_vmat(0,3)(40),
			mult_vmat(0,4)(40),
			mult_vmat(1,3)(40),
			mult_vmat(1,1)(41)
		);

		mult_vmat(1,4)(40) <= mult_vmat(0,5)(40);
		mult_vmat(1,5)(40) <= mult_vmat(0,6)(40);
		mult_vmat(1,6)(40) <= mult_vmat(0,7)(40);
		mult_vmat(1,7)(40) <= mult_vmat(0,8)(40);
		mult_vmat(1,8)(40) <= mult_vmat(0,9)(40);
		mult_vmat(1,9)(40) <= mult_vmat(0,10)(40);
		mult_vmat(1,10)(40) <= mult_vmat(0,11)(40);
		mult_vmat(1,11)(40) <= mult_vmat(0,12)(40);
		mult_vmat(1,12)(40) <= mult_vmat(0,13)(40);

		-- COLUMN 42

		FA_0_41_1: FA PORT MAP (
			mult_vmat(0,0)(41),
			mult_vmat(0,1)(41),
			mult_vmat(0,2)(41),
			mult_vmat(1,2)(41),
			mult_vmat(1,0)(42)
		);

		mult_vmat(1,3)(41) <= mult_vmat(0,3)(41);
		mult_vmat(1,4)(41) <= mult_vmat(0,4)(41);
		mult_vmat(1,5)(41) <= mult_vmat(0,5)(41);
		mult_vmat(1,6)(41) <= mult_vmat(0,6)(41);
		mult_vmat(1,7)(41) <= mult_vmat(0,7)(41);
		mult_vmat(1,8)(41) <= mult_vmat(0,8)(41);
		mult_vmat(1,9)(41) <= mult_vmat(0,9)(41);
		mult_vmat(1,10)(41) <= mult_vmat(0,10)(41);
		mult_vmat(1,11)(41) <= mult_vmat(0,11)(41);
		mult_vmat(1,12)(41) <= mult_vmat(0,12)(41);

		-- COLUMN 43

		HA_0_42: HA PORT MAP (
			mult_vmat(0,0)(42),
			mult_vmat(0,1)(42),
			mult_vmat(1,1)(42),
			mult_vmat(1,0)(43)
		);

		mult_vmat(1,2)(42) <= mult_vmat(0,2)(42);
		mult_vmat(1,3)(42) <= mult_vmat(0,3)(42);
		mult_vmat(1,4)(42) <= mult_vmat(0,4)(42);
		mult_vmat(1,5)(42) <= mult_vmat(0,5)(42);
		mult_vmat(1,6)(42) <= mult_vmat(0,6)(42);
		mult_vmat(1,7)(42) <= mult_vmat(0,7)(42);
		mult_vmat(1,8)(42) <= mult_vmat(0,8)(42);
		mult_vmat(1,9)(42) <= mult_vmat(0,9)(42);
		mult_vmat(1,10)(42) <= mult_vmat(0,10)(42);
		mult_vmat(1,11)(42) <= mult_vmat(0,11)(42);
		mult_vmat(1,12)(42) <= mult_vmat(0,12)(42);

		-- COLUMN 44
		mult_vmat(1,1)(43) <= mult_vmat(0,0)(43);
		mult_vmat(1,2)(43) <= mult_vmat(0,1)(43);
		mult_vmat(1,3)(43) <= mult_vmat(0,2)(43);
		mult_vmat(1,4)(43) <= mult_vmat(0,3)(43);
		mult_vmat(1,5)(43) <= mult_vmat(0,4)(43);
		mult_vmat(1,6)(43) <= mult_vmat(0,5)(43);
		mult_vmat(1,7)(43) <= mult_vmat(0,6)(43);
		mult_vmat(1,8)(43) <= mult_vmat(0,7)(43);
		mult_vmat(1,9)(43) <= mult_vmat(0,8)(43);
		mult_vmat(1,10)(43) <= mult_vmat(0,9)(43);
		mult_vmat(1,11)(43) <= mult_vmat(0,10)(43);
		mult_vmat(1,12)(43) <= mult_vmat(0,11)(43);

		-- COLUMN 45
		mult_vmat(1,0)(44) <= mult_vmat(0,0)(44);
		mult_vmat(1,1)(44) <= mult_vmat(0,1)(44);
		mult_vmat(1,2)(44) <= mult_vmat(0,2)(44);
		mult_vmat(1,3)(44) <= mult_vmat(0,3)(44);
		mult_vmat(1,4)(44) <= mult_vmat(0,4)(44);
		mult_vmat(1,5)(44) <= mult_vmat(0,5)(44);
		mult_vmat(1,6)(44) <= mult_vmat(0,6)(44);
		mult_vmat(1,7)(44) <= mult_vmat(0,7)(44);
		mult_vmat(1,8)(44) <= mult_vmat(0,8)(44);
		mult_vmat(1,9)(44) <= mult_vmat(0,9)(44);
		mult_vmat(1,10)(44) <= mult_vmat(0,10)(44);
		mult_vmat(1,11)(44) <= mult_vmat(0,11)(44);

		-- COLUMN 46
		mult_vmat(1,0)(45) <= mult_vmat(0,0)(45);
		mult_vmat(1,1)(45) <= mult_vmat(0,1)(45);
		mult_vmat(1,2)(45) <= mult_vmat(0,2)(45);
		mult_vmat(1,3)(45) <= mult_vmat(0,3)(45);
		mult_vmat(1,4)(45) <= mult_vmat(0,4)(45);
		mult_vmat(1,5)(45) <= mult_vmat(0,5)(45);
		mult_vmat(1,6)(45) <= mult_vmat(0,6)(45);
		mult_vmat(1,7)(45) <= mult_vmat(0,7)(45);
		mult_vmat(1,8)(45) <= mult_vmat(0,8)(45);
		mult_vmat(1,9)(45) <= mult_vmat(0,9)(45);
		mult_vmat(1,10)(45) <= mult_vmat(0,10)(45);

		-- COLUMN 47
		mult_vmat(1,0)(46) <= mult_vmat(0,0)(46);
		mult_vmat(1,1)(46) <= mult_vmat(0,1)(46);
		mult_vmat(1,2)(46) <= mult_vmat(0,2)(46);
		mult_vmat(1,3)(46) <= mult_vmat(0,3)(46);
		mult_vmat(1,4)(46) <= mult_vmat(0,4)(46);
		mult_vmat(1,5)(46) <= mult_vmat(0,5)(46);
		mult_vmat(1,6)(46) <= mult_vmat(0,6)(46);
		mult_vmat(1,7)(46) <= mult_vmat(0,7)(46);
		mult_vmat(1,8)(46) <= mult_vmat(0,8)(46);
		mult_vmat(1,9)(46) <= mult_vmat(0,9)(46);
		mult_vmat(1,10)(46) <= mult_vmat(0,10)(46);

		-- COLUMN 48
		mult_vmat(1,0)(47) <= mult_vmat(0,0)(47);
		mult_vmat(1,1)(47) <= mult_vmat(0,1)(47);
		mult_vmat(1,2)(47) <= mult_vmat(0,2)(47);
		mult_vmat(1,3)(47) <= mult_vmat(0,3)(47);
		mult_vmat(1,4)(47) <= mult_vmat(0,4)(47);
		mult_vmat(1,5)(47) <= mult_vmat(0,5)(47);
		mult_vmat(1,6)(47) <= mult_vmat(0,6)(47);
		mult_vmat(1,7)(47) <= mult_vmat(0,7)(47);
		mult_vmat(1,8)(47) <= mult_vmat(0,8)(47);
		mult_vmat(1,9)(47) <= mult_vmat(0,9)(47);

		-- COLUMN 49
		mult_vmat(1,0)(48) <= mult_vmat(0,0)(48);
		mult_vmat(1,1)(48) <= mult_vmat(0,1)(48);
		mult_vmat(1,2)(48) <= mult_vmat(0,2)(48);
		mult_vmat(1,3)(48) <= mult_vmat(0,3)(48);
		mult_vmat(1,4)(48) <= mult_vmat(0,4)(48);
		mult_vmat(1,5)(48) <= mult_vmat(0,5)(48);
		mult_vmat(1,6)(48) <= mult_vmat(0,6)(48);
		mult_vmat(1,7)(48) <= mult_vmat(0,7)(48);
		mult_vmat(1,8)(48) <= mult_vmat(0,8)(48);
		mult_vmat(1,9)(48) <= mult_vmat(0,9)(48);

		-- COLUMN 50
		mult_vmat(1,0)(49) <= mult_vmat(0,0)(49);
		mult_vmat(1,1)(49) <= mult_vmat(0,1)(49);
		mult_vmat(1,2)(49) <= mult_vmat(0,2)(49);
		mult_vmat(1,3)(49) <= mult_vmat(0,3)(49);
		mult_vmat(1,4)(49) <= mult_vmat(0,4)(49);
		mult_vmat(1,5)(49) <= mult_vmat(0,5)(49);
		mult_vmat(1,6)(49) <= mult_vmat(0,6)(49);
		mult_vmat(1,7)(49) <= mult_vmat(0,7)(49);
		mult_vmat(1,8)(49) <= mult_vmat(0,8)(49);

		-- COLUMN 51
		mult_vmat(1,0)(50) <= mult_vmat(0,0)(50);
		mult_vmat(1,1)(50) <= mult_vmat(0,1)(50);
		mult_vmat(1,2)(50) <= mult_vmat(0,2)(50);
		mult_vmat(1,3)(50) <= mult_vmat(0,3)(50);
		mult_vmat(1,4)(50) <= mult_vmat(0,4)(50);
		mult_vmat(1,5)(50) <= mult_vmat(0,5)(50);
		mult_vmat(1,6)(50) <= mult_vmat(0,6)(50);
		mult_vmat(1,7)(50) <= mult_vmat(0,7)(50);
		mult_vmat(1,8)(50) <= mult_vmat(0,8)(50);

		-- COLUMN 52
		mult_vmat(1,0)(51) <= mult_vmat(0,0)(51);
		mult_vmat(1,1)(51) <= mult_vmat(0,1)(51);
		mult_vmat(1,2)(51) <= mult_vmat(0,2)(51);
		mult_vmat(1,3)(51) <= mult_vmat(0,3)(51);
		mult_vmat(1,4)(51) <= mult_vmat(0,4)(51);
		mult_vmat(1,5)(51) <= mult_vmat(0,5)(51);
		mult_vmat(1,6)(51) <= mult_vmat(0,6)(51);
		mult_vmat(1,7)(51) <= mult_vmat(0,7)(51);

		-- COLUMN 53
		mult_vmat(1,0)(52) <= mult_vmat(0,0)(52);
		mult_vmat(1,1)(52) <= mult_vmat(0,1)(52);
		mult_vmat(1,2)(52) <= mult_vmat(0,2)(52);
		mult_vmat(1,3)(52) <= mult_vmat(0,3)(52);
		mult_vmat(1,4)(52) <= mult_vmat(0,4)(52);
		mult_vmat(1,5)(52) <= mult_vmat(0,5)(52);
		mult_vmat(1,6)(52) <= mult_vmat(0,6)(52);
		mult_vmat(1,7)(52) <= mult_vmat(0,7)(52);

		-- COLUMN 54
		mult_vmat(1,0)(53) <= mult_vmat(0,0)(53);
		mult_vmat(1,1)(53) <= mult_vmat(0,1)(53);
		mult_vmat(1,2)(53) <= mult_vmat(0,2)(53);
		mult_vmat(1,3)(53) <= mult_vmat(0,3)(53);
		mult_vmat(1,4)(53) <= mult_vmat(0,4)(53);
		mult_vmat(1,5)(53) <= mult_vmat(0,5)(53);
		mult_vmat(1,6)(53) <= mult_vmat(0,6)(53);

		-- COLUMN 55
		mult_vmat(1,0)(54) <= mult_vmat(0,0)(54);
		mult_vmat(1,1)(54) <= mult_vmat(0,1)(54);
		mult_vmat(1,2)(54) <= mult_vmat(0,2)(54);
		mult_vmat(1,3)(54) <= mult_vmat(0,3)(54);
		mult_vmat(1,4)(54) <= mult_vmat(0,4)(54);
		mult_vmat(1,5)(54) <= mult_vmat(0,5)(54);
		mult_vmat(1,6)(54) <= mult_vmat(0,6)(54);

		-- COLUMN 56
		mult_vmat(1,0)(55) <= mult_vmat(0,0)(55);
		mult_vmat(1,1)(55) <= mult_vmat(0,1)(55);
		mult_vmat(1,2)(55) <= mult_vmat(0,2)(55);
		mult_vmat(1,3)(55) <= mult_vmat(0,3)(55);
		mult_vmat(1,4)(55) <= mult_vmat(0,4)(55);
		mult_vmat(1,5)(55) <= mult_vmat(0,5)(55);

		-- COLUMN 57
		mult_vmat(1,0)(56) <= mult_vmat(0,0)(56);
		mult_vmat(1,1)(56) <= mult_vmat(0,1)(56);
		mult_vmat(1,2)(56) <= mult_vmat(0,2)(56);
		mult_vmat(1,3)(56) <= mult_vmat(0,3)(56);
		mult_vmat(1,4)(56) <= mult_vmat(0,4)(56);
		mult_vmat(1,5)(56) <= mult_vmat(0,5)(56);

		-- COLUMN 58
		mult_vmat(1,0)(57) <= mult_vmat(0,0)(57);
		mult_vmat(1,1)(57) <= mult_vmat(0,1)(57);
		mult_vmat(1,2)(57) <= mult_vmat(0,2)(57);
		mult_vmat(1,3)(57) <= mult_vmat(0,3)(57);
		mult_vmat(1,4)(57) <= mult_vmat(0,4)(57);

		-- COLUMN 59
		mult_vmat(1,0)(58) <= mult_vmat(0,0)(58);
		mult_vmat(1,1)(58) <= mult_vmat(0,1)(58);
		mult_vmat(1,2)(58) <= mult_vmat(0,2)(58);
		mult_vmat(1,3)(58) <= mult_vmat(0,3)(58);
		mult_vmat(1,4)(58) <= mult_vmat(0,4)(58);

		-- COLUMN 60
		mult_vmat(1,0)(59) <= mult_vmat(0,0)(59);
		mult_vmat(1,1)(59) <= mult_vmat(0,1)(59);
		mult_vmat(1,2)(59) <= mult_vmat(0,2)(59);
		mult_vmat(1,3)(59) <= mult_vmat(0,3)(59);

		-- COLUMN 61
		mult_vmat(1,0)(60) <= mult_vmat(0,0)(60);
		mult_vmat(1,1)(60) <= mult_vmat(0,1)(60);
		mult_vmat(1,2)(60) <= mult_vmat(0,2)(60);
		mult_vmat(1,3)(60) <= mult_vmat(0,3)(60);

		-- COLUMN 62
		mult_vmat(1,0)(61) <= mult_vmat(0,0)(61);
		mult_vmat(1,1)(61) <= mult_vmat(0,1)(61);
		mult_vmat(1,2)(61) <= mult_vmat(0,2)(61);

		-- COLUMN 63
		mult_vmat(1,0)(62) <= mult_vmat(0,0)(62);
		mult_vmat(1,1)(62) <= mult_vmat(0,1)(62);
		mult_vmat(1,2)(62) <= mult_vmat(0,2)(62);

		-- COLUMN 64
		mult_vmat(1,0)(63) <= mult_vmat(0,0)(63);
		mult_vmat(1,1)(63) <= mult_vmat(0,1)(63);


	------------------------------------------
	-- LEVEL 2
	------------------------------------------


		-- COLUMN 1
		mult_vmat(2,0)(0) <= mult_vmat(1,0)(0);
		mult_vmat(2,1)(0) <= mult_vmat(1,1)(0);

		-- COLUMN 2
		mult_vmat(2,0)(1) <= mult_vmat(1,0)(1);

		-- COLUMN 3
		mult_vmat(2,0)(2) <= mult_vmat(1,0)(2);
		mult_vmat(2,1)(2) <= mult_vmat(1,1)(2);
		mult_vmat(2,2)(2) <= mult_vmat(1,2)(2);

		-- COLUMN 4
		mult_vmat(2,0)(3) <= mult_vmat(1,0)(3);
		mult_vmat(2,1)(3) <= mult_vmat(1,1)(3);

		-- COLUMN 5
		mult_vmat(2,0)(4) <= mult_vmat(1,0)(4);
		mult_vmat(2,1)(4) <= mult_vmat(1,1)(4);
		mult_vmat(2,2)(4) <= mult_vmat(1,2)(4);
		mult_vmat(2,3)(4) <= mult_vmat(1,3)(4);

		-- COLUMN 6
		mult_vmat(2,0)(5) <= mult_vmat(1,0)(5);
		mult_vmat(2,1)(5) <= mult_vmat(1,1)(5);
		mult_vmat(2,2)(5) <= mult_vmat(1,2)(5);

		-- COLUMN 7
		mult_vmat(2,0)(6) <= mult_vmat(1,0)(6);
		mult_vmat(2,1)(6) <= mult_vmat(1,1)(6);
		mult_vmat(2,2)(6) <= mult_vmat(1,2)(6);
		mult_vmat(2,3)(6) <= mult_vmat(1,3)(6);
		mult_vmat(2,4)(6) <= mult_vmat(1,4)(6);

		-- COLUMN 8
		mult_vmat(2,0)(7) <= mult_vmat(1,0)(7);
		mult_vmat(2,1)(7) <= mult_vmat(1,1)(7);
		mult_vmat(2,2)(7) <= mult_vmat(1,2)(7);
		mult_vmat(2,3)(7) <= mult_vmat(1,3)(7);

		-- COLUMN 9
		mult_vmat(2,0)(8) <= mult_vmat(1,0)(8);
		mult_vmat(2,1)(8) <= mult_vmat(1,1)(8);
		mult_vmat(2,2)(8) <= mult_vmat(1,2)(8);
		mult_vmat(2,3)(8) <= mult_vmat(1,3)(8);
		mult_vmat(2,4)(8) <= mult_vmat(1,4)(8);
		mult_vmat(2,5)(8) <= mult_vmat(1,5)(8);

		-- COLUMN 10
		mult_vmat(2,0)(9) <= mult_vmat(1,0)(9);
		mult_vmat(2,1)(9) <= mult_vmat(1,1)(9);
		mult_vmat(2,2)(9) <= mult_vmat(1,2)(9);
		mult_vmat(2,3)(9) <= mult_vmat(1,3)(9);
		mult_vmat(2,4)(9) <= mult_vmat(1,4)(9);

		-- COLUMN 11
		mult_vmat(2,0)(10) <= mult_vmat(1,0)(10);
		mult_vmat(2,1)(10) <= mult_vmat(1,1)(10);
		mult_vmat(2,2)(10) <= mult_vmat(1,2)(10);
		mult_vmat(2,3)(10) <= mult_vmat(1,3)(10);
		mult_vmat(2,4)(10) <= mult_vmat(1,4)(10);
		mult_vmat(2,5)(10) <= mult_vmat(1,5)(10);
		mult_vmat(2,6)(10) <= mult_vmat(1,6)(10);

		-- COLUMN 12
		mult_vmat(2,0)(11) <= mult_vmat(1,0)(11);
		mult_vmat(2,1)(11) <= mult_vmat(1,1)(11);
		mult_vmat(2,2)(11) <= mult_vmat(1,2)(11);
		mult_vmat(2,3)(11) <= mult_vmat(1,3)(11);
		mult_vmat(2,4)(11) <= mult_vmat(1,4)(11);
		mult_vmat(2,5)(11) <= mult_vmat(1,5)(11);

		-- COLUMN 13
		mult_vmat(2,0)(12) <= mult_vmat(1,0)(12);
		mult_vmat(2,1)(12) <= mult_vmat(1,1)(12);
		mult_vmat(2,2)(12) <= mult_vmat(1,2)(12);
		mult_vmat(2,3)(12) <= mult_vmat(1,3)(12);
		mult_vmat(2,4)(12) <= mult_vmat(1,4)(12);
		mult_vmat(2,5)(12) <= mult_vmat(1,5)(12);
		mult_vmat(2,6)(12) <= mult_vmat(1,6)(12);
		mult_vmat(2,7)(12) <= mult_vmat(1,7)(12);

		-- COLUMN 14
		mult_vmat(2,0)(13) <= mult_vmat(1,0)(13);
		mult_vmat(2,1)(13) <= mult_vmat(1,1)(13);
		mult_vmat(2,2)(13) <= mult_vmat(1,2)(13);
		mult_vmat(2,3)(13) <= mult_vmat(1,3)(13);
		mult_vmat(2,4)(13) <= mult_vmat(1,4)(13);
		mult_vmat(2,5)(13) <= mult_vmat(1,5)(13);
		mult_vmat(2,6)(13) <= mult_vmat(1,6)(13);

		-- COLUMN 15
		mult_vmat(2,0)(14) <= mult_vmat(1,0)(14);
		mult_vmat(2,1)(14) <= mult_vmat(1,1)(14);
		mult_vmat(2,2)(14) <= mult_vmat(1,2)(14);
		mult_vmat(2,3)(14) <= mult_vmat(1,3)(14);
		mult_vmat(2,4)(14) <= mult_vmat(1,4)(14);
		mult_vmat(2,5)(14) <= mult_vmat(1,5)(14);
		mult_vmat(2,6)(14) <= mult_vmat(1,6)(14);
		mult_vmat(2,7)(14) <= mult_vmat(1,7)(14);
		mult_vmat(2,8)(14) <= mult_vmat(1,8)(14);

		-- COLUMN 16
		mult_vmat(2,0)(15) <= mult_vmat(1,0)(15);
		mult_vmat(2,1)(15) <= mult_vmat(1,1)(15);
		mult_vmat(2,2)(15) <= mult_vmat(1,2)(15);
		mult_vmat(2,3)(15) <= mult_vmat(1,3)(15);
		mult_vmat(2,4)(15) <= mult_vmat(1,4)(15);
		mult_vmat(2,5)(15) <= mult_vmat(1,5)(15);
		mult_vmat(2,6)(15) <= mult_vmat(1,6)(15);
		mult_vmat(2,7)(15) <= mult_vmat(1,7)(15);

		-- COLUMN 17

		HA_1_16: HA PORT MAP (
			mult_vmat(1,0)(16),
			mult_vmat(1,1)(16),
			mult_vmat(2,0)(16),
			mult_vmat(2,0)(17)
		);

		mult_vmat(2,1)(16) <= mult_vmat(1,2)(16);
		mult_vmat(2,2)(16) <= mult_vmat(1,3)(16);
		mult_vmat(2,3)(16) <= mult_vmat(1,4)(16);
		mult_vmat(2,4)(16) <= mult_vmat(1,5)(16);
		mult_vmat(2,5)(16) <= mult_vmat(1,6)(16);
		mult_vmat(2,6)(16) <= mult_vmat(1,7)(16);
		mult_vmat(2,7)(16) <= mult_vmat(1,8)(16);
		mult_vmat(2,8)(16) <= mult_vmat(1,9)(16);

		-- COLUMN 18

		HA_1_17: HA PORT MAP (
			mult_vmat(1,0)(17),
			mult_vmat(1,1)(17),
			mult_vmat(2,1)(17),
			mult_vmat(2,0)(18)
		);

		mult_vmat(2,2)(17) <= mult_vmat(1,2)(17);
		mult_vmat(2,3)(17) <= mult_vmat(1,3)(17);
		mult_vmat(2,4)(17) <= mult_vmat(1,4)(17);
		mult_vmat(2,5)(17) <= mult_vmat(1,5)(17);
		mult_vmat(2,6)(17) <= mult_vmat(1,6)(17);
		mult_vmat(2,7)(17) <= mult_vmat(1,7)(17);
		mult_vmat(2,8)(17) <= mult_vmat(1,8)(17);

		-- COLUMN 19

		FA_1_18_1: FA PORT MAP (
			mult_vmat(1,0)(18),
			mult_vmat(1,1)(18),
			mult_vmat(1,2)(18),
			mult_vmat(2,1)(18),
			mult_vmat(2,0)(19)
		);


		HA_1_18: HA PORT MAP (
			mult_vmat(1,3)(18),
			mult_vmat(1,4)(18),
			mult_vmat(2,2)(18),
			mult_vmat(2,1)(19)
		);

		mult_vmat(2,3)(18) <= mult_vmat(1,5)(18);
		mult_vmat(2,4)(18) <= mult_vmat(1,6)(18);
		mult_vmat(2,5)(18) <= mult_vmat(1,7)(18);
		mult_vmat(2,6)(18) <= mult_vmat(1,8)(18);
		mult_vmat(2,7)(18) <= mult_vmat(1,9)(18);
		mult_vmat(2,8)(18) <= mult_vmat(1,10)(18);

		-- COLUMN 20

		FA_1_19_1: FA PORT MAP (
			mult_vmat(1,0)(19),
			mult_vmat(1,1)(19),
			mult_vmat(1,2)(19),
			mult_vmat(2,2)(19),
			mult_vmat(2,0)(20)
		);


		HA_1_19: HA PORT MAP (
			mult_vmat(1,3)(19),
			mult_vmat(1,4)(19),
			mult_vmat(2,3)(19),
			mult_vmat(2,1)(20)
		);

		mult_vmat(2,4)(19) <= mult_vmat(1,5)(19);
		mult_vmat(2,5)(19) <= mult_vmat(1,6)(19);
		mult_vmat(2,6)(19) <= mult_vmat(1,7)(19);
		mult_vmat(2,7)(19) <= mult_vmat(1,8)(19);
		mult_vmat(2,8)(19) <= mult_vmat(1,9)(19);

		-- COLUMN 21

		FA_1_20_1: FA PORT MAP (
			mult_vmat(1,0)(20),
			mult_vmat(1,1)(20),
			mult_vmat(1,2)(20),
			mult_vmat(2,2)(20),
			mult_vmat(2,0)(21)
		);


		FA_1_20_2: FA PORT MAP (
			mult_vmat(1,3)(20),
			mult_vmat(1,4)(20),
			mult_vmat(1,5)(20),
			mult_vmat(2,3)(20),
			mult_vmat(2,1)(21)
		);


		HA_1_20: HA PORT MAP (
			mult_vmat(1,6)(20),
			mult_vmat(1,7)(20),
			mult_vmat(2,4)(20),
			mult_vmat(2,2)(21)
		);

		mult_vmat(2,5)(20) <= mult_vmat(1,8)(20);
		mult_vmat(2,6)(20) <= mult_vmat(1,9)(20);
		mult_vmat(2,7)(20) <= mult_vmat(1,10)(20);
		mult_vmat(2,8)(20) <= mult_vmat(1,11)(20);

		-- COLUMN 22

		FA_1_21_1: FA PORT MAP (
			mult_vmat(1,0)(21),
			mult_vmat(1,1)(21),
			mult_vmat(1,2)(21),
			mult_vmat(2,3)(21),
			mult_vmat(2,0)(22)
		);


		FA_1_21_2: FA PORT MAP (
			mult_vmat(1,3)(21),
			mult_vmat(1,4)(21),
			mult_vmat(1,5)(21),
			mult_vmat(2,4)(21),
			mult_vmat(2,1)(22)
		);


		HA_1_21: HA PORT MAP (
			mult_vmat(1,6)(21),
			mult_vmat(1,7)(21),
			mult_vmat(2,5)(21),
			mult_vmat(2,2)(22)
		);

		mult_vmat(2,6)(21) <= mult_vmat(1,8)(21);
		mult_vmat(2,7)(21) <= mult_vmat(1,9)(21);
		mult_vmat(2,8)(21) <= mult_vmat(1,10)(21);

		-- COLUMN 23

		FA_1_22_1: FA PORT MAP (
			mult_vmat(1,0)(22),
			mult_vmat(1,1)(22),
			mult_vmat(1,2)(22),
			mult_vmat(2,3)(22),
			mult_vmat(2,0)(23)
		);


		FA_1_22_2: FA PORT MAP (
			mult_vmat(1,3)(22),
			mult_vmat(1,4)(22),
			mult_vmat(1,5)(22),
			mult_vmat(2,4)(22),
			mult_vmat(2,1)(23)
		);


		FA_1_22_3: FA PORT MAP (
			mult_vmat(1,6)(22),
			mult_vmat(1,7)(22),
			mult_vmat(1,8)(22),
			mult_vmat(2,5)(22),
			mult_vmat(2,2)(23)
		);


		HA_1_22: HA PORT MAP (
			mult_vmat(1,9)(22),
			mult_vmat(1,10)(22),
			mult_vmat(2,6)(22),
			mult_vmat(2,3)(23)
		);

		mult_vmat(2,7)(22) <= mult_vmat(1,11)(22);
		mult_vmat(2,8)(22) <= mult_vmat(1,12)(22);

		-- COLUMN 24

		FA_1_23_1: FA PORT MAP (
			mult_vmat(1,0)(23),
			mult_vmat(1,1)(23),
			mult_vmat(1,2)(23),
			mult_vmat(2,4)(23),
			mult_vmat(2,0)(24)
		);


		FA_1_23_2: FA PORT MAP (
			mult_vmat(1,3)(23),
			mult_vmat(1,4)(23),
			mult_vmat(1,5)(23),
			mult_vmat(2,5)(23),
			mult_vmat(2,1)(24)
		);


		FA_1_23_3: FA PORT MAP (
			mult_vmat(1,6)(23),
			mult_vmat(1,7)(23),
			mult_vmat(1,8)(23),
			mult_vmat(2,6)(23),
			mult_vmat(2,2)(24)
		);


		HA_1_23: HA PORT MAP (
			mult_vmat(1,9)(23),
			mult_vmat(1,10)(23),
			mult_vmat(2,7)(23),
			mult_vmat(2,3)(24)
		);

		mult_vmat(2,8)(23) <= mult_vmat(1,11)(23);

		-- COLUMN 25

		FA_1_24_1: FA PORT MAP (
			mult_vmat(1,0)(24),
			mult_vmat(1,1)(24),
			mult_vmat(1,2)(24),
			mult_vmat(2,4)(24),
			mult_vmat(2,0)(25)
		);


		FA_1_24_2: FA PORT MAP (
			mult_vmat(1,3)(24),
			mult_vmat(1,4)(24),
			mult_vmat(1,5)(24),
			mult_vmat(2,5)(24),
			mult_vmat(2,1)(25)
		);


		FA_1_24_3: FA PORT MAP (
			mult_vmat(1,6)(24),
			mult_vmat(1,7)(24),
			mult_vmat(1,8)(24),
			mult_vmat(2,6)(24),
			mult_vmat(2,2)(25)
		);


		FA_1_24_4: FA PORT MAP (
			mult_vmat(1,9)(24),
			mult_vmat(1,10)(24),
			mult_vmat(1,11)(24),
			mult_vmat(2,7)(24),
			mult_vmat(2,3)(25)
		);

		mult_vmat(2,8)(24) <= mult_vmat(1,12)(24);

		-- COLUMN 26

		FA_1_25_1: FA PORT MAP (
			mult_vmat(1,0)(25),
			mult_vmat(1,1)(25),
			mult_vmat(1,2)(25),
			mult_vmat(2,4)(25),
			mult_vmat(2,0)(26)
		);


		FA_1_25_2: FA PORT MAP (
			mult_vmat(1,3)(25),
			mult_vmat(1,4)(25),
			mult_vmat(1,5)(25),
			mult_vmat(2,5)(25),
			mult_vmat(2,1)(26)
		);


		FA_1_25_3: FA PORT MAP (
			mult_vmat(1,6)(25),
			mult_vmat(1,7)(25),
			mult_vmat(1,8)(25),
			mult_vmat(2,6)(25),
			mult_vmat(2,2)(26)
		);


		FA_1_25_4: FA PORT MAP (
			mult_vmat(1,9)(25),
			mult_vmat(1,10)(25),
			mult_vmat(1,11)(25),
			mult_vmat(2,7)(25),
			mult_vmat(2,3)(26)
		);

		mult_vmat(2,8)(25) <= mult_vmat(1,12)(25);

		-- COLUMN 27

		FA_1_26_1: FA PORT MAP (
			mult_vmat(1,0)(26),
			mult_vmat(1,1)(26),
			mult_vmat(1,2)(26),
			mult_vmat(2,4)(26),
			mult_vmat(2,0)(27)
		);


		FA_1_26_2: FA PORT MAP (
			mult_vmat(1,3)(26),
			mult_vmat(1,4)(26),
			mult_vmat(1,5)(26),
			mult_vmat(2,5)(26),
			mult_vmat(2,1)(27)
		);


		FA_1_26_3: FA PORT MAP (
			mult_vmat(1,6)(26),
			mult_vmat(1,7)(26),
			mult_vmat(1,8)(26),
			mult_vmat(2,6)(26),
			mult_vmat(2,2)(27)
		);


		FA_1_26_4: FA PORT MAP (
			mult_vmat(1,9)(26),
			mult_vmat(1,10)(26),
			mult_vmat(1,11)(26),
			mult_vmat(2,7)(26),
			mult_vmat(2,3)(27)
		);

		mult_vmat(2,8)(26) <= mult_vmat(1,12)(26);

		-- COLUMN 28

		FA_1_27_1: FA PORT MAP (
			mult_vmat(1,0)(27),
			mult_vmat(1,1)(27),
			mult_vmat(1,2)(27),
			mult_vmat(2,4)(27),
			mult_vmat(2,0)(28)
		);


		FA_1_27_2: FA PORT MAP (
			mult_vmat(1,3)(27),
			mult_vmat(1,4)(27),
			mult_vmat(1,5)(27),
			mult_vmat(2,5)(27),
			mult_vmat(2,1)(28)
		);


		FA_1_27_3: FA PORT MAP (
			mult_vmat(1,6)(27),
			mult_vmat(1,7)(27),
			mult_vmat(1,8)(27),
			mult_vmat(2,6)(27),
			mult_vmat(2,2)(28)
		);


		FA_1_27_4: FA PORT MAP (
			mult_vmat(1,9)(27),
			mult_vmat(1,10)(27),
			mult_vmat(1,11)(27),
			mult_vmat(2,7)(27),
			mult_vmat(2,3)(28)
		);

		mult_vmat(2,8)(27) <= mult_vmat(1,12)(27);

		-- COLUMN 29

		FA_1_28_1: FA PORT MAP (
			mult_vmat(1,0)(28),
			mult_vmat(1,1)(28),
			mult_vmat(1,2)(28),
			mult_vmat(2,4)(28),
			mult_vmat(2,0)(29)
		);


		FA_1_28_2: FA PORT MAP (
			mult_vmat(1,3)(28),
			mult_vmat(1,4)(28),
			mult_vmat(1,5)(28),
			mult_vmat(2,5)(28),
			mult_vmat(2,1)(29)
		);


		FA_1_28_3: FA PORT MAP (
			mult_vmat(1,6)(28),
			mult_vmat(1,7)(28),
			mult_vmat(1,8)(28),
			mult_vmat(2,6)(28),
			mult_vmat(2,2)(29)
		);


		FA_1_28_4: FA PORT MAP (
			mult_vmat(1,9)(28),
			mult_vmat(1,10)(28),
			mult_vmat(1,11)(28),
			mult_vmat(2,7)(28),
			mult_vmat(2,3)(29)
		);

		mult_vmat(2,8)(28) <= mult_vmat(1,12)(28);

		-- COLUMN 30

		FA_1_29_1: FA PORT MAP (
			mult_vmat(1,0)(29),
			mult_vmat(1,1)(29),
			mult_vmat(1,2)(29),
			mult_vmat(2,4)(29),
			mult_vmat(2,0)(30)
		);


		FA_1_29_2: FA PORT MAP (
			mult_vmat(1,3)(29),
			mult_vmat(1,4)(29),
			mult_vmat(1,5)(29),
			mult_vmat(2,5)(29),
			mult_vmat(2,1)(30)
		);


		FA_1_29_3: FA PORT MAP (
			mult_vmat(1,6)(29),
			mult_vmat(1,7)(29),
			mult_vmat(1,8)(29),
			mult_vmat(2,6)(29),
			mult_vmat(2,2)(30)
		);


		FA_1_29_4: FA PORT MAP (
			mult_vmat(1,9)(29),
			mult_vmat(1,10)(29),
			mult_vmat(1,11)(29),
			mult_vmat(2,7)(29),
			mult_vmat(2,3)(30)
		);

		mult_vmat(2,8)(29) <= mult_vmat(1,12)(29);

		-- COLUMN 31

		FA_1_30_1: FA PORT MAP (
			mult_vmat(1,0)(30),
			mult_vmat(1,1)(30),
			mult_vmat(1,2)(30),
			mult_vmat(2,4)(30),
			mult_vmat(2,0)(31)
		);


		FA_1_30_2: FA PORT MAP (
			mult_vmat(1,3)(30),
			mult_vmat(1,4)(30),
			mult_vmat(1,5)(30),
			mult_vmat(2,5)(30),
			mult_vmat(2,1)(31)
		);


		FA_1_30_3: FA PORT MAP (
			mult_vmat(1,6)(30),
			mult_vmat(1,7)(30),
			mult_vmat(1,8)(30),
			mult_vmat(2,6)(30),
			mult_vmat(2,2)(31)
		);


		FA_1_30_4: FA PORT MAP (
			mult_vmat(1,9)(30),
			mult_vmat(1,10)(30),
			mult_vmat(1,11)(30),
			mult_vmat(2,7)(30),
			mult_vmat(2,3)(31)
		);

		mult_vmat(2,8)(30) <= mult_vmat(1,12)(30);

		-- COLUMN 32

		FA_1_31_1: FA PORT MAP (
			mult_vmat(1,0)(31),
			mult_vmat(1,1)(31),
			mult_vmat(1,2)(31),
			mult_vmat(2,4)(31),
			mult_vmat(2,0)(32)
		);


		FA_1_31_2: FA PORT MAP (
			mult_vmat(1,3)(31),
			mult_vmat(1,4)(31),
			mult_vmat(1,5)(31),
			mult_vmat(2,5)(31),
			mult_vmat(2,1)(32)
		);


		FA_1_31_3: FA PORT MAP (
			mult_vmat(1,6)(31),
			mult_vmat(1,7)(31),
			mult_vmat(1,8)(31),
			mult_vmat(2,6)(31),
			mult_vmat(2,2)(32)
		);


		FA_1_31_4: FA PORT MAP (
			mult_vmat(1,9)(31),
			mult_vmat(1,10)(31),
			mult_vmat(1,11)(31),
			mult_vmat(2,7)(31),
			mult_vmat(2,3)(32)
		);

		mult_vmat(2,8)(31) <= mult_vmat(1,12)(31);

		-- COLUMN 33

		FA_1_32_1: FA PORT MAP (
			mult_vmat(1,0)(32),
			mult_vmat(1,1)(32),
			mult_vmat(1,2)(32),
			mult_vmat(2,4)(32),
			mult_vmat(2,0)(33)
		);


		FA_1_32_2: FA PORT MAP (
			mult_vmat(1,3)(32),
			mult_vmat(1,4)(32),
			mult_vmat(1,5)(32),
			mult_vmat(2,5)(32),
			mult_vmat(2,1)(33)
		);


		FA_1_32_3: FA PORT MAP (
			mult_vmat(1,6)(32),
			mult_vmat(1,7)(32),
			mult_vmat(1,8)(32),
			mult_vmat(2,6)(32),
			mult_vmat(2,2)(33)
		);


		FA_1_32_4: FA PORT MAP (
			mult_vmat(1,9)(32),
			mult_vmat(1,10)(32),
			mult_vmat(1,11)(32),
			mult_vmat(2,7)(32),
			mult_vmat(2,3)(33)
		);

		mult_vmat(2,8)(32) <= mult_vmat(1,12)(32);

		-- COLUMN 34

		FA_1_33_1: FA PORT MAP (
			mult_vmat(1,0)(33),
			mult_vmat(1,1)(33),
			mult_vmat(1,2)(33),
			mult_vmat(2,4)(33),
			mult_vmat(2,0)(34)
		);


		FA_1_33_2: FA PORT MAP (
			mult_vmat(1,3)(33),
			mult_vmat(1,4)(33),
			mult_vmat(1,5)(33),
			mult_vmat(2,5)(33),
			mult_vmat(2,1)(34)
		);


		FA_1_33_3: FA PORT MAP (
			mult_vmat(1,6)(33),
			mult_vmat(1,7)(33),
			mult_vmat(1,8)(33),
			mult_vmat(2,6)(33),
			mult_vmat(2,2)(34)
		);


		FA_1_33_4: FA PORT MAP (
			mult_vmat(1,9)(33),
			mult_vmat(1,10)(33),
			mult_vmat(1,11)(33),
			mult_vmat(2,7)(33),
			mult_vmat(2,3)(34)
		);

		mult_vmat(2,8)(33) <= mult_vmat(1,12)(33);

		-- COLUMN 35

		FA_1_34_1: FA PORT MAP (
			mult_vmat(1,0)(34),
			mult_vmat(1,1)(34),
			mult_vmat(1,2)(34),
			mult_vmat(2,4)(34),
			mult_vmat(2,0)(35)
		);


		FA_1_34_2: FA PORT MAP (
			mult_vmat(1,3)(34),
			mult_vmat(1,4)(34),
			mult_vmat(1,5)(34),
			mult_vmat(2,5)(34),
			mult_vmat(2,1)(35)
		);


		FA_1_34_3: FA PORT MAP (
			mult_vmat(1,6)(34),
			mult_vmat(1,7)(34),
			mult_vmat(1,8)(34),
			mult_vmat(2,6)(34),
			mult_vmat(2,2)(35)
		);


		FA_1_34_4: FA PORT MAP (
			mult_vmat(1,9)(34),
			mult_vmat(1,10)(34),
			mult_vmat(1,11)(34),
			mult_vmat(2,7)(34),
			mult_vmat(2,3)(35)
		);

		mult_vmat(2,8)(34) <= mult_vmat(1,12)(34);

		-- COLUMN 36

		FA_1_35_1: FA PORT MAP (
			mult_vmat(1,0)(35),
			mult_vmat(1,1)(35),
			mult_vmat(1,2)(35),
			mult_vmat(2,4)(35),
			mult_vmat(2,0)(36)
		);


		FA_1_35_2: FA PORT MAP (
			mult_vmat(1,3)(35),
			mult_vmat(1,4)(35),
			mult_vmat(1,5)(35),
			mult_vmat(2,5)(35),
			mult_vmat(2,1)(36)
		);


		FA_1_35_3: FA PORT MAP (
			mult_vmat(1,6)(35),
			mult_vmat(1,7)(35),
			mult_vmat(1,8)(35),
			mult_vmat(2,6)(35),
			mult_vmat(2,2)(36)
		);


		FA_1_35_4: FA PORT MAP (
			mult_vmat(1,9)(35),
			mult_vmat(1,10)(35),
			mult_vmat(1,11)(35),
			mult_vmat(2,7)(35),
			mult_vmat(2,3)(36)
		);

		mult_vmat(2,8)(35) <= mult_vmat(1,12)(35);

		-- COLUMN 37

		FA_1_36_1: FA PORT MAP (
			mult_vmat(1,0)(36),
			mult_vmat(1,1)(36),
			mult_vmat(1,2)(36),
			mult_vmat(2,4)(36),
			mult_vmat(2,0)(37)
		);


		FA_1_36_2: FA PORT MAP (
			mult_vmat(1,3)(36),
			mult_vmat(1,4)(36),
			mult_vmat(1,5)(36),
			mult_vmat(2,5)(36),
			mult_vmat(2,1)(37)
		);


		FA_1_36_3: FA PORT MAP (
			mult_vmat(1,6)(36),
			mult_vmat(1,7)(36),
			mult_vmat(1,8)(36),
			mult_vmat(2,6)(36),
			mult_vmat(2,2)(37)
		);


		FA_1_36_4: FA PORT MAP (
			mult_vmat(1,9)(36),
			mult_vmat(1,10)(36),
			mult_vmat(1,11)(36),
			mult_vmat(2,7)(36),
			mult_vmat(2,3)(37)
		);

		mult_vmat(2,8)(36) <= mult_vmat(1,12)(36);

		-- COLUMN 38

		FA_1_37_1: FA PORT MAP (
			mult_vmat(1,0)(37),
			mult_vmat(1,1)(37),
			mult_vmat(1,2)(37),
			mult_vmat(2,4)(37),
			mult_vmat(2,0)(38)
		);


		FA_1_37_2: FA PORT MAP (
			mult_vmat(1,3)(37),
			mult_vmat(1,4)(37),
			mult_vmat(1,5)(37),
			mult_vmat(2,5)(37),
			mult_vmat(2,1)(38)
		);


		FA_1_37_3: FA PORT MAP (
			mult_vmat(1,6)(37),
			mult_vmat(1,7)(37),
			mult_vmat(1,8)(37),
			mult_vmat(2,6)(37),
			mult_vmat(2,2)(38)
		);


		FA_1_37_4: FA PORT MAP (
			mult_vmat(1,9)(37),
			mult_vmat(1,10)(37),
			mult_vmat(1,11)(37),
			mult_vmat(2,7)(37),
			mult_vmat(2,3)(38)
		);

		mult_vmat(2,8)(37) <= mult_vmat(1,12)(37);

		-- COLUMN 39

		FA_1_38_1: FA PORT MAP (
			mult_vmat(1,0)(38),
			mult_vmat(1,1)(38),
			mult_vmat(1,2)(38),
			mult_vmat(2,4)(38),
			mult_vmat(2,0)(39)
		);


		FA_1_38_2: FA PORT MAP (
			mult_vmat(1,3)(38),
			mult_vmat(1,4)(38),
			mult_vmat(1,5)(38),
			mult_vmat(2,5)(38),
			mult_vmat(2,1)(39)
		);


		FA_1_38_3: FA PORT MAP (
			mult_vmat(1,6)(38),
			mult_vmat(1,7)(38),
			mult_vmat(1,8)(38),
			mult_vmat(2,6)(38),
			mult_vmat(2,2)(39)
		);


		FA_1_38_4: FA PORT MAP (
			mult_vmat(1,9)(38),
			mult_vmat(1,10)(38),
			mult_vmat(1,11)(38),
			mult_vmat(2,7)(38),
			mult_vmat(2,3)(39)
		);

		mult_vmat(2,8)(38) <= mult_vmat(1,12)(38);

		-- COLUMN 40

		FA_1_39_1: FA PORT MAP (
			mult_vmat(1,0)(39),
			mult_vmat(1,1)(39),
			mult_vmat(1,2)(39),
			mult_vmat(2,4)(39),
			mult_vmat(2,0)(40)
		);


		FA_1_39_2: FA PORT MAP (
			mult_vmat(1,3)(39),
			mult_vmat(1,4)(39),
			mult_vmat(1,5)(39),
			mult_vmat(2,5)(39),
			mult_vmat(2,1)(40)
		);


		FA_1_39_3: FA PORT MAP (
			mult_vmat(1,6)(39),
			mult_vmat(1,7)(39),
			mult_vmat(1,8)(39),
			mult_vmat(2,6)(39),
			mult_vmat(2,2)(40)
		);


		FA_1_39_4: FA PORT MAP (
			mult_vmat(1,9)(39),
			mult_vmat(1,10)(39),
			mult_vmat(1,11)(39),
			mult_vmat(2,7)(39),
			mult_vmat(2,3)(40)
		);

		mult_vmat(2,8)(39) <= mult_vmat(1,12)(39);

		-- COLUMN 41

		FA_1_40_1: FA PORT MAP (
			mult_vmat(1,0)(40),
			mult_vmat(1,1)(40),
			mult_vmat(1,2)(40),
			mult_vmat(2,4)(40),
			mult_vmat(2,0)(41)
		);


		FA_1_40_2: FA PORT MAP (
			mult_vmat(1,3)(40),
			mult_vmat(1,4)(40),
			mult_vmat(1,5)(40),
			mult_vmat(2,5)(40),
			mult_vmat(2,1)(41)
		);


		FA_1_40_3: FA PORT MAP (
			mult_vmat(1,6)(40),
			mult_vmat(1,7)(40),
			mult_vmat(1,8)(40),
			mult_vmat(2,6)(40),
			mult_vmat(2,2)(41)
		);


		FA_1_40_4: FA PORT MAP (
			mult_vmat(1,9)(40),
			mult_vmat(1,10)(40),
			mult_vmat(1,11)(40),
			mult_vmat(2,7)(40),
			mult_vmat(2,3)(41)
		);

		mult_vmat(2,8)(40) <= mult_vmat(1,12)(40);

		-- COLUMN 42

		FA_1_41_1: FA PORT MAP (
			mult_vmat(1,0)(41),
			mult_vmat(1,1)(41),
			mult_vmat(1,2)(41),
			mult_vmat(2,4)(41),
			mult_vmat(2,0)(42)
		);


		FA_1_41_2: FA PORT MAP (
			mult_vmat(1,3)(41),
			mult_vmat(1,4)(41),
			mult_vmat(1,5)(41),
			mult_vmat(2,5)(41),
			mult_vmat(2,1)(42)
		);


		FA_1_41_3: FA PORT MAP (
			mult_vmat(1,6)(41),
			mult_vmat(1,7)(41),
			mult_vmat(1,8)(41),
			mult_vmat(2,6)(41),
			mult_vmat(2,2)(42)
		);


		FA_1_41_4: FA PORT MAP (
			mult_vmat(1,9)(41),
			mult_vmat(1,10)(41),
			mult_vmat(1,11)(41),
			mult_vmat(2,7)(41),
			mult_vmat(2,3)(42)
		);

		mult_vmat(2,8)(41) <= mult_vmat(1,12)(41);

		-- COLUMN 43

		FA_1_42_1: FA PORT MAP (
			mult_vmat(1,0)(42),
			mult_vmat(1,1)(42),
			mult_vmat(1,2)(42),
			mult_vmat(2,4)(42),
			mult_vmat(2,0)(43)
		);


		FA_1_42_2: FA PORT MAP (
			mult_vmat(1,3)(42),
			mult_vmat(1,4)(42),
			mult_vmat(1,5)(42),
			mult_vmat(2,5)(42),
			mult_vmat(2,1)(43)
		);


		FA_1_42_3: FA PORT MAP (
			mult_vmat(1,6)(42),
			mult_vmat(1,7)(42),
			mult_vmat(1,8)(42),
			mult_vmat(2,6)(42),
			mult_vmat(2,2)(43)
		);


		FA_1_42_4: FA PORT MAP (
			mult_vmat(1,9)(42),
			mult_vmat(1,10)(42),
			mult_vmat(1,11)(42),
			mult_vmat(2,7)(42),
			mult_vmat(2,3)(43)
		);

		mult_vmat(2,8)(42) <= mult_vmat(1,12)(42);

		-- COLUMN 44

		FA_1_43_1: FA PORT MAP (
			mult_vmat(1,0)(43),
			mult_vmat(1,1)(43),
			mult_vmat(1,2)(43),
			mult_vmat(2,4)(43),
			mult_vmat(2,0)(44)
		);


		FA_1_43_2: FA PORT MAP (
			mult_vmat(1,3)(43),
			mult_vmat(1,4)(43),
			mult_vmat(1,5)(43),
			mult_vmat(2,5)(43),
			mult_vmat(2,1)(44)
		);


		FA_1_43_3: FA PORT MAP (
			mult_vmat(1,6)(43),
			mult_vmat(1,7)(43),
			mult_vmat(1,8)(43),
			mult_vmat(2,6)(43),
			mult_vmat(2,2)(44)
		);


		FA_1_43_4: FA PORT MAP (
			mult_vmat(1,9)(43),
			mult_vmat(1,10)(43),
			mult_vmat(1,11)(43),
			mult_vmat(2,7)(43),
			mult_vmat(2,3)(44)
		);

		mult_vmat(2,8)(43) <= mult_vmat(1,12)(43);

		-- COLUMN 45

		FA_1_44_1: FA PORT MAP (
			mult_vmat(1,0)(44),
			mult_vmat(1,1)(44),
			mult_vmat(1,2)(44),
			mult_vmat(2,4)(44),
			mult_vmat(2,0)(45)
		);


		FA_1_44_2: FA PORT MAP (
			mult_vmat(1,3)(44),
			mult_vmat(1,4)(44),
			mult_vmat(1,5)(44),
			mult_vmat(2,5)(44),
			mult_vmat(2,1)(45)
		);


		FA_1_44_3: FA PORT MAP (
			mult_vmat(1,6)(44),
			mult_vmat(1,7)(44),
			mult_vmat(1,8)(44),
			mult_vmat(2,6)(44),
			mult_vmat(2,2)(45)
		);


		HA_1_44: HA PORT MAP (
			mult_vmat(1,9)(44),
			mult_vmat(1,10)(44),
			mult_vmat(2,7)(44),
			mult_vmat(2,3)(45)
		);

		mult_vmat(2,8)(44) <= mult_vmat(1,11)(44);

		-- COLUMN 46

		FA_1_45_1: FA PORT MAP (
			mult_vmat(1,0)(45),
			mult_vmat(1,1)(45),
			mult_vmat(1,2)(45),
			mult_vmat(2,4)(45),
			mult_vmat(2,0)(46)
		);


		FA_1_45_2: FA PORT MAP (
			mult_vmat(1,3)(45),
			mult_vmat(1,4)(45),
			mult_vmat(1,5)(45),
			mult_vmat(2,5)(45),
			mult_vmat(2,1)(46)
		);


		FA_1_45_3: FA PORT MAP (
			mult_vmat(1,6)(45),
			mult_vmat(1,7)(45),
			mult_vmat(1,8)(45),
			mult_vmat(2,6)(45),
			mult_vmat(2,2)(46)
		);

		mult_vmat(2,7)(45) <= mult_vmat(1,9)(45);
		mult_vmat(2,8)(45) <= mult_vmat(1,10)(45);

		-- COLUMN 47

		FA_1_46_1: FA PORT MAP (
			mult_vmat(1,0)(46),
			mult_vmat(1,1)(46),
			mult_vmat(1,2)(46),
			mult_vmat(2,3)(46),
			mult_vmat(2,0)(47)
		);


		FA_1_46_2: FA PORT MAP (
			mult_vmat(1,3)(46),
			mult_vmat(1,4)(46),
			mult_vmat(1,5)(46),
			mult_vmat(2,4)(46),
			mult_vmat(2,1)(47)
		);


		HA_1_46: HA PORT MAP (
			mult_vmat(1,6)(46),
			mult_vmat(1,7)(46),
			mult_vmat(2,5)(46),
			mult_vmat(2,2)(47)
		);

		mult_vmat(2,6)(46) <= mult_vmat(1,8)(46);
		mult_vmat(2,7)(46) <= mult_vmat(1,9)(46);
		mult_vmat(2,8)(46) <= mult_vmat(1,10)(46);

		-- COLUMN 48

		FA_1_47_1: FA PORT MAP (
			mult_vmat(1,0)(47),
			mult_vmat(1,1)(47),
			mult_vmat(1,2)(47),
			mult_vmat(2,3)(47),
			mult_vmat(2,0)(48)
		);


		FA_1_47_2: FA PORT MAP (
			mult_vmat(1,3)(47),
			mult_vmat(1,4)(47),
			mult_vmat(1,5)(47),
			mult_vmat(2,4)(47),
			mult_vmat(2,1)(48)
		);

		mult_vmat(2,5)(47) <= mult_vmat(1,6)(47);
		mult_vmat(2,6)(47) <= mult_vmat(1,7)(47);
		mult_vmat(2,7)(47) <= mult_vmat(1,8)(47);
		mult_vmat(2,8)(47) <= mult_vmat(1,9)(47);

		-- COLUMN 49

		FA_1_48_1: FA PORT MAP (
			mult_vmat(1,0)(48),
			mult_vmat(1,1)(48),
			mult_vmat(1,2)(48),
			mult_vmat(2,2)(48),
			mult_vmat(2,0)(49)
		);


		HA_1_48: HA PORT MAP (
			mult_vmat(1,3)(48),
			mult_vmat(1,4)(48),
			mult_vmat(2,3)(48),
			mult_vmat(2,1)(49)
		);

		mult_vmat(2,4)(48) <= mult_vmat(1,5)(48);
		mult_vmat(2,5)(48) <= mult_vmat(1,6)(48);
		mult_vmat(2,6)(48) <= mult_vmat(1,7)(48);
		mult_vmat(2,7)(48) <= mult_vmat(1,8)(48);
		mult_vmat(2,8)(48) <= mult_vmat(1,9)(48);

		-- COLUMN 50

		FA_1_49_1: FA PORT MAP (
			mult_vmat(1,0)(49),
			mult_vmat(1,1)(49),
			mult_vmat(1,2)(49),
			mult_vmat(2,2)(49),
			mult_vmat(2,0)(50)
		);

		mult_vmat(2,3)(49) <= mult_vmat(1,3)(49);
		mult_vmat(2,4)(49) <= mult_vmat(1,4)(49);
		mult_vmat(2,5)(49) <= mult_vmat(1,5)(49);
		mult_vmat(2,6)(49) <= mult_vmat(1,6)(49);
		mult_vmat(2,7)(49) <= mult_vmat(1,7)(49);
		mult_vmat(2,8)(49) <= mult_vmat(1,8)(49);

		-- COLUMN 51

		HA_1_50: HA PORT MAP (
			mult_vmat(1,0)(50),
			mult_vmat(1,1)(50),
			mult_vmat(2,1)(50),
			mult_vmat(2,0)(51)
		);

		mult_vmat(2,2)(50) <= mult_vmat(1,2)(50);
		mult_vmat(2,3)(50) <= mult_vmat(1,3)(50);
		mult_vmat(2,4)(50) <= mult_vmat(1,4)(50);
		mult_vmat(2,5)(50) <= mult_vmat(1,5)(50);
		mult_vmat(2,6)(50) <= mult_vmat(1,6)(50);
		mult_vmat(2,7)(50) <= mult_vmat(1,7)(50);
		mult_vmat(2,8)(50) <= mult_vmat(1,8)(50);

		-- COLUMN 52
		mult_vmat(2,1)(51) <= mult_vmat(1,0)(51);
		mult_vmat(2,2)(51) <= mult_vmat(1,1)(51);
		mult_vmat(2,3)(51) <= mult_vmat(1,2)(51);
		mult_vmat(2,4)(51) <= mult_vmat(1,3)(51);
		mult_vmat(2,5)(51) <= mult_vmat(1,4)(51);
		mult_vmat(2,6)(51) <= mult_vmat(1,5)(51);
		mult_vmat(2,7)(51) <= mult_vmat(1,6)(51);
		mult_vmat(2,8)(51) <= mult_vmat(1,7)(51);

		-- COLUMN 53
		mult_vmat(2,0)(52) <= mult_vmat(1,0)(52);
		mult_vmat(2,1)(52) <= mult_vmat(1,1)(52);
		mult_vmat(2,2)(52) <= mult_vmat(1,2)(52);
		mult_vmat(2,3)(52) <= mult_vmat(1,3)(52);
		mult_vmat(2,4)(52) <= mult_vmat(1,4)(52);
		mult_vmat(2,5)(52) <= mult_vmat(1,5)(52);
		mult_vmat(2,6)(52) <= mult_vmat(1,6)(52);
		mult_vmat(2,7)(52) <= mult_vmat(1,7)(52);

		-- COLUMN 54
		mult_vmat(2,0)(53) <= mult_vmat(1,0)(53);
		mult_vmat(2,1)(53) <= mult_vmat(1,1)(53);
		mult_vmat(2,2)(53) <= mult_vmat(1,2)(53);
		mult_vmat(2,3)(53) <= mult_vmat(1,3)(53);
		mult_vmat(2,4)(53) <= mult_vmat(1,4)(53);
		mult_vmat(2,5)(53) <= mult_vmat(1,5)(53);
		mult_vmat(2,6)(53) <= mult_vmat(1,6)(53);

		-- COLUMN 55
		mult_vmat(2,0)(54) <= mult_vmat(1,0)(54);
		mult_vmat(2,1)(54) <= mult_vmat(1,1)(54);
		mult_vmat(2,2)(54) <= mult_vmat(1,2)(54);
		mult_vmat(2,3)(54) <= mult_vmat(1,3)(54);
		mult_vmat(2,4)(54) <= mult_vmat(1,4)(54);
		mult_vmat(2,5)(54) <= mult_vmat(1,5)(54);
		mult_vmat(2,6)(54) <= mult_vmat(1,6)(54);

		-- COLUMN 56
		mult_vmat(2,0)(55) <= mult_vmat(1,0)(55);
		mult_vmat(2,1)(55) <= mult_vmat(1,1)(55);
		mult_vmat(2,2)(55) <= mult_vmat(1,2)(55);
		mult_vmat(2,3)(55) <= mult_vmat(1,3)(55);
		mult_vmat(2,4)(55) <= mult_vmat(1,4)(55);
		mult_vmat(2,5)(55) <= mult_vmat(1,5)(55);

		-- COLUMN 57
		mult_vmat(2,0)(56) <= mult_vmat(1,0)(56);
		mult_vmat(2,1)(56) <= mult_vmat(1,1)(56);
		mult_vmat(2,2)(56) <= mult_vmat(1,2)(56);
		mult_vmat(2,3)(56) <= mult_vmat(1,3)(56);
		mult_vmat(2,4)(56) <= mult_vmat(1,4)(56);
		mult_vmat(2,5)(56) <= mult_vmat(1,5)(56);

		-- COLUMN 58
		mult_vmat(2,0)(57) <= mult_vmat(1,0)(57);
		mult_vmat(2,1)(57) <= mult_vmat(1,1)(57);
		mult_vmat(2,2)(57) <= mult_vmat(1,2)(57);
		mult_vmat(2,3)(57) <= mult_vmat(1,3)(57);
		mult_vmat(2,4)(57) <= mult_vmat(1,4)(57);

		-- COLUMN 59
		mult_vmat(2,0)(58) <= mult_vmat(1,0)(58);
		mult_vmat(2,1)(58) <= mult_vmat(1,1)(58);
		mult_vmat(2,2)(58) <= mult_vmat(1,2)(58);
		mult_vmat(2,3)(58) <= mult_vmat(1,3)(58);
		mult_vmat(2,4)(58) <= mult_vmat(1,4)(58);

		-- COLUMN 60
		mult_vmat(2,0)(59) <= mult_vmat(1,0)(59);
		mult_vmat(2,1)(59) <= mult_vmat(1,1)(59);
		mult_vmat(2,2)(59) <= mult_vmat(1,2)(59);
		mult_vmat(2,3)(59) <= mult_vmat(1,3)(59);

		-- COLUMN 61
		mult_vmat(2,0)(60) <= mult_vmat(1,0)(60);
		mult_vmat(2,1)(60) <= mult_vmat(1,1)(60);
		mult_vmat(2,2)(60) <= mult_vmat(1,2)(60);
		mult_vmat(2,3)(60) <= mult_vmat(1,3)(60);

		-- COLUMN 62
		mult_vmat(2,0)(61) <= mult_vmat(1,0)(61);
		mult_vmat(2,1)(61) <= mult_vmat(1,1)(61);
		mult_vmat(2,2)(61) <= mult_vmat(1,2)(61);

		-- COLUMN 63
		mult_vmat(2,0)(62) <= mult_vmat(1,0)(62);
		mult_vmat(2,1)(62) <= mult_vmat(1,1)(62);
		mult_vmat(2,2)(62) <= mult_vmat(1,2)(62);

		-- COLUMN 64
		mult_vmat(2,0)(63) <= mult_vmat(1,0)(63);
		mult_vmat(2,1)(63) <= mult_vmat(1,1)(63);


	------------------------------------------
	-- LEVEL 3
	------------------------------------------


		-- COLUMN 1
		mult_vmat(3,0)(0) <= mult_vmat(2,0)(0);
		mult_vmat(3,1)(0) <= mult_vmat(2,1)(0);

		-- COLUMN 2
		mult_vmat(3,0)(1) <= mult_vmat(2,0)(1);

		-- COLUMN 3
		mult_vmat(3,0)(2) <= mult_vmat(2,0)(2);
		mult_vmat(3,1)(2) <= mult_vmat(2,1)(2);
		mult_vmat(3,2)(2) <= mult_vmat(2,2)(2);

		-- COLUMN 4
		mult_vmat(3,0)(3) <= mult_vmat(2,0)(3);
		mult_vmat(3,1)(3) <= mult_vmat(2,1)(3);

		-- COLUMN 5
		mult_vmat(3,0)(4) <= mult_vmat(2,0)(4);
		mult_vmat(3,1)(4) <= mult_vmat(2,1)(4);
		mult_vmat(3,2)(4) <= mult_vmat(2,2)(4);
		mult_vmat(3,3)(4) <= mult_vmat(2,3)(4);

		-- COLUMN 6
		mult_vmat(3,0)(5) <= mult_vmat(2,0)(5);
		mult_vmat(3,1)(5) <= mult_vmat(2,1)(5);
		mult_vmat(3,2)(5) <= mult_vmat(2,2)(5);

		-- COLUMN 7
		mult_vmat(3,0)(6) <= mult_vmat(2,0)(6);
		mult_vmat(3,1)(6) <= mult_vmat(2,1)(6);
		mult_vmat(3,2)(6) <= mult_vmat(2,2)(6);
		mult_vmat(3,3)(6) <= mult_vmat(2,3)(6);
		mult_vmat(3,4)(6) <= mult_vmat(2,4)(6);

		-- COLUMN 8
		mult_vmat(3,0)(7) <= mult_vmat(2,0)(7);
		mult_vmat(3,1)(7) <= mult_vmat(2,1)(7);
		mult_vmat(3,2)(7) <= mult_vmat(2,2)(7);
		mult_vmat(3,3)(7) <= mult_vmat(2,3)(7);

		-- COLUMN 9
		mult_vmat(3,0)(8) <= mult_vmat(2,0)(8);
		mult_vmat(3,1)(8) <= mult_vmat(2,1)(8);
		mult_vmat(3,2)(8) <= mult_vmat(2,2)(8);
		mult_vmat(3,3)(8) <= mult_vmat(2,3)(8);
		mult_vmat(3,4)(8) <= mult_vmat(2,4)(8);
		mult_vmat(3,5)(8) <= mult_vmat(2,5)(8);

		-- COLUMN 10
		mult_vmat(3,0)(9) <= mult_vmat(2,0)(9);
		mult_vmat(3,1)(9) <= mult_vmat(2,1)(9);
		mult_vmat(3,2)(9) <= mult_vmat(2,2)(9);
		mult_vmat(3,3)(9) <= mult_vmat(2,3)(9);
		mult_vmat(3,4)(9) <= mult_vmat(2,4)(9);

		-- COLUMN 11

		HA_2_10: HA PORT MAP (
			mult_vmat(2,0)(10),
			mult_vmat(2,1)(10),
			mult_vmat(3,0)(10),
			mult_vmat(3,0)(11)
		);

		mult_vmat(3,1)(10) <= mult_vmat(2,2)(10);
		mult_vmat(3,2)(10) <= mult_vmat(2,3)(10);
		mult_vmat(3,3)(10) <= mult_vmat(2,4)(10);
		mult_vmat(3,4)(10) <= mult_vmat(2,5)(10);
		mult_vmat(3,5)(10) <= mult_vmat(2,6)(10);

		-- COLUMN 12

		HA_2_11: HA PORT MAP (
			mult_vmat(2,0)(11),
			mult_vmat(2,1)(11),
			mult_vmat(3,1)(11),
			mult_vmat(3,0)(12)
		);

		mult_vmat(3,2)(11) <= mult_vmat(2,2)(11);
		mult_vmat(3,3)(11) <= mult_vmat(2,3)(11);
		mult_vmat(3,4)(11) <= mult_vmat(2,4)(11);
		mult_vmat(3,5)(11) <= mult_vmat(2,5)(11);

		-- COLUMN 13

		FA_2_12_1: FA PORT MAP (
			mult_vmat(2,0)(12),
			mult_vmat(2,1)(12),
			mult_vmat(2,2)(12),
			mult_vmat(3,1)(12),
			mult_vmat(3,0)(13)
		);


		HA_2_12: HA PORT MAP (
			mult_vmat(2,3)(12),
			mult_vmat(2,4)(12),
			mult_vmat(3,2)(12),
			mult_vmat(3,1)(13)
		);

		mult_vmat(3,3)(12) <= mult_vmat(2,5)(12);
		mult_vmat(3,4)(12) <= mult_vmat(2,6)(12);
		mult_vmat(3,5)(12) <= mult_vmat(2,7)(12);

		-- COLUMN 14

		FA_2_13_1: FA PORT MAP (
			mult_vmat(2,0)(13),
			mult_vmat(2,1)(13),
			mult_vmat(2,2)(13),
			mult_vmat(3,2)(13),
			mult_vmat(3,0)(14)
		);


		HA_2_13: HA PORT MAP (
			mult_vmat(2,3)(13),
			mult_vmat(2,4)(13),
			mult_vmat(3,3)(13),
			mult_vmat(3,1)(14)
		);

		mult_vmat(3,4)(13) <= mult_vmat(2,5)(13);
		mult_vmat(3,5)(13) <= mult_vmat(2,6)(13);

		-- COLUMN 15

		FA_2_14_1: FA PORT MAP (
			mult_vmat(2,0)(14),
			mult_vmat(2,1)(14),
			mult_vmat(2,2)(14),
			mult_vmat(3,2)(14),
			mult_vmat(3,0)(15)
		);


		FA_2_14_2: FA PORT MAP (
			mult_vmat(2,3)(14),
			mult_vmat(2,4)(14),
			mult_vmat(2,5)(14),
			mult_vmat(3,3)(14),
			mult_vmat(3,1)(15)
		);


		HA_2_14: HA PORT MAP (
			mult_vmat(2,6)(14),
			mult_vmat(2,7)(14),
			mult_vmat(3,4)(14),
			mult_vmat(3,2)(15)
		);

		mult_vmat(3,5)(14) <= mult_vmat(2,8)(14);

		-- COLUMN 16

		FA_2_15_1: FA PORT MAP (
			mult_vmat(2,0)(15),
			mult_vmat(2,1)(15),
			mult_vmat(2,2)(15),
			mult_vmat(3,3)(15),
			mult_vmat(3,0)(16)
		);


		FA_2_15_2: FA PORT MAP (
			mult_vmat(2,3)(15),
			mult_vmat(2,4)(15),
			mult_vmat(2,5)(15),
			mult_vmat(3,4)(15),
			mult_vmat(3,1)(16)
		);


		HA_2_15: HA PORT MAP (
			mult_vmat(2,6)(15),
			mult_vmat(2,7)(15),
			mult_vmat(3,5)(15),
			mult_vmat(3,2)(16)
		);


		-- COLUMN 17

		FA_2_16_1: FA PORT MAP (
			mult_vmat(2,0)(16),
			mult_vmat(2,1)(16),
			mult_vmat(2,2)(16),
			mult_vmat(3,3)(16),
			mult_vmat(3,0)(17)
		);


		FA_2_16_2: FA PORT MAP (
			mult_vmat(2,3)(16),
			mult_vmat(2,4)(16),
			mult_vmat(2,5)(16),
			mult_vmat(3,4)(16),
			mult_vmat(3,1)(17)
		);


		FA_2_16_3: FA PORT MAP (
			mult_vmat(2,6)(16),
			mult_vmat(2,7)(16),
			mult_vmat(2,8)(16),
			mult_vmat(3,5)(16),
			mult_vmat(3,2)(17)
		);


		-- COLUMN 18

		FA_2_17_1: FA PORT MAP (
			mult_vmat(2,0)(17),
			mult_vmat(2,1)(17),
			mult_vmat(2,2)(17),
			mult_vmat(3,3)(17),
			mult_vmat(3,0)(18)
		);


		FA_2_17_2: FA PORT MAP (
			mult_vmat(2,3)(17),
			mult_vmat(2,4)(17),
			mult_vmat(2,5)(17),
			mult_vmat(3,4)(17),
			mult_vmat(3,1)(18)
		);


		FA_2_17_3: FA PORT MAP (
			mult_vmat(2,6)(17),
			mult_vmat(2,7)(17),
			mult_vmat(2,8)(17),
			mult_vmat(3,5)(17),
			mult_vmat(3,2)(18)
		);


		-- COLUMN 19

		FA_2_18_1: FA PORT MAP (
			mult_vmat(2,0)(18),
			mult_vmat(2,1)(18),
			mult_vmat(2,2)(18),
			mult_vmat(3,3)(18),
			mult_vmat(3,0)(19)
		);


		FA_2_18_2: FA PORT MAP (
			mult_vmat(2,3)(18),
			mult_vmat(2,4)(18),
			mult_vmat(2,5)(18),
			mult_vmat(3,4)(18),
			mult_vmat(3,1)(19)
		);


		FA_2_18_3: FA PORT MAP (
			mult_vmat(2,6)(18),
			mult_vmat(2,7)(18),
			mult_vmat(2,8)(18),
			mult_vmat(3,5)(18),
			mult_vmat(3,2)(19)
		);


		-- COLUMN 20

		FA_2_19_1: FA PORT MAP (
			mult_vmat(2,0)(19),
			mult_vmat(2,1)(19),
			mult_vmat(2,2)(19),
			mult_vmat(3,3)(19),
			mult_vmat(3,0)(20)
		);


		FA_2_19_2: FA PORT MAP (
			mult_vmat(2,3)(19),
			mult_vmat(2,4)(19),
			mult_vmat(2,5)(19),
			mult_vmat(3,4)(19),
			mult_vmat(3,1)(20)
		);


		FA_2_19_3: FA PORT MAP (
			mult_vmat(2,6)(19),
			mult_vmat(2,7)(19),
			mult_vmat(2,8)(19),
			mult_vmat(3,5)(19),
			mult_vmat(3,2)(20)
		);


		-- COLUMN 21

		FA_2_20_1: FA PORT MAP (
			mult_vmat(2,0)(20),
			mult_vmat(2,1)(20),
			mult_vmat(2,2)(20),
			mult_vmat(3,3)(20),
			mult_vmat(3,0)(21)
		);


		FA_2_20_2: FA PORT MAP (
			mult_vmat(2,3)(20),
			mult_vmat(2,4)(20),
			mult_vmat(2,5)(20),
			mult_vmat(3,4)(20),
			mult_vmat(3,1)(21)
		);


		FA_2_20_3: FA PORT MAP (
			mult_vmat(2,6)(20),
			mult_vmat(2,7)(20),
			mult_vmat(2,8)(20),
			mult_vmat(3,5)(20),
			mult_vmat(3,2)(21)
		);


		-- COLUMN 22

		FA_2_21_1: FA PORT MAP (
			mult_vmat(2,0)(21),
			mult_vmat(2,1)(21),
			mult_vmat(2,2)(21),
			mult_vmat(3,3)(21),
			mult_vmat(3,0)(22)
		);


		FA_2_21_2: FA PORT MAP (
			mult_vmat(2,3)(21),
			mult_vmat(2,4)(21),
			mult_vmat(2,5)(21),
			mult_vmat(3,4)(21),
			mult_vmat(3,1)(22)
		);


		FA_2_21_3: FA PORT MAP (
			mult_vmat(2,6)(21),
			mult_vmat(2,7)(21),
			mult_vmat(2,8)(21),
			mult_vmat(3,5)(21),
			mult_vmat(3,2)(22)
		);


		-- COLUMN 23

		FA_2_22_1: FA PORT MAP (
			mult_vmat(2,0)(22),
			mult_vmat(2,1)(22),
			mult_vmat(2,2)(22),
			mult_vmat(3,3)(22),
			mult_vmat(3,0)(23)
		);


		FA_2_22_2: FA PORT MAP (
			mult_vmat(2,3)(22),
			mult_vmat(2,4)(22),
			mult_vmat(2,5)(22),
			mult_vmat(3,4)(22),
			mult_vmat(3,1)(23)
		);


		FA_2_22_3: FA PORT MAP (
			mult_vmat(2,6)(22),
			mult_vmat(2,7)(22),
			mult_vmat(2,8)(22),
			mult_vmat(3,5)(22),
			mult_vmat(3,2)(23)
		);


		-- COLUMN 24

		FA_2_23_1: FA PORT MAP (
			mult_vmat(2,0)(23),
			mult_vmat(2,1)(23),
			mult_vmat(2,2)(23),
			mult_vmat(3,3)(23),
			mult_vmat(3,0)(24)
		);


		FA_2_23_2: FA PORT MAP (
			mult_vmat(2,3)(23),
			mult_vmat(2,4)(23),
			mult_vmat(2,5)(23),
			mult_vmat(3,4)(23),
			mult_vmat(3,1)(24)
		);


		FA_2_23_3: FA PORT MAP (
			mult_vmat(2,6)(23),
			mult_vmat(2,7)(23),
			mult_vmat(2,8)(23),
			mult_vmat(3,5)(23),
			mult_vmat(3,2)(24)
		);


		-- COLUMN 25

		FA_2_24_1: FA PORT MAP (
			mult_vmat(2,0)(24),
			mult_vmat(2,1)(24),
			mult_vmat(2,2)(24),
			mult_vmat(3,3)(24),
			mult_vmat(3,0)(25)
		);


		FA_2_24_2: FA PORT MAP (
			mult_vmat(2,3)(24),
			mult_vmat(2,4)(24),
			mult_vmat(2,5)(24),
			mult_vmat(3,4)(24),
			mult_vmat(3,1)(25)
		);


		FA_2_24_3: FA PORT MAP (
			mult_vmat(2,6)(24),
			mult_vmat(2,7)(24),
			mult_vmat(2,8)(24),
			mult_vmat(3,5)(24),
			mult_vmat(3,2)(25)
		);


		-- COLUMN 26

		FA_2_25_1: FA PORT MAP (
			mult_vmat(2,0)(25),
			mult_vmat(2,1)(25),
			mult_vmat(2,2)(25),
			mult_vmat(3,3)(25),
			mult_vmat(3,0)(26)
		);


		FA_2_25_2: FA PORT MAP (
			mult_vmat(2,3)(25),
			mult_vmat(2,4)(25),
			mult_vmat(2,5)(25),
			mult_vmat(3,4)(25),
			mult_vmat(3,1)(26)
		);


		FA_2_25_3: FA PORT MAP (
			mult_vmat(2,6)(25),
			mult_vmat(2,7)(25),
			mult_vmat(2,8)(25),
			mult_vmat(3,5)(25),
			mult_vmat(3,2)(26)
		);


		-- COLUMN 27

		FA_2_26_1: FA PORT MAP (
			mult_vmat(2,0)(26),
			mult_vmat(2,1)(26),
			mult_vmat(2,2)(26),
			mult_vmat(3,3)(26),
			mult_vmat(3,0)(27)
		);


		FA_2_26_2: FA PORT MAP (
			mult_vmat(2,3)(26),
			mult_vmat(2,4)(26),
			mult_vmat(2,5)(26),
			mult_vmat(3,4)(26),
			mult_vmat(3,1)(27)
		);


		FA_2_26_3: FA PORT MAP (
			mult_vmat(2,6)(26),
			mult_vmat(2,7)(26),
			mult_vmat(2,8)(26),
			mult_vmat(3,5)(26),
			mult_vmat(3,2)(27)
		);


		-- COLUMN 28

		FA_2_27_1: FA PORT MAP (
			mult_vmat(2,0)(27),
			mult_vmat(2,1)(27),
			mult_vmat(2,2)(27),
			mult_vmat(3,3)(27),
			mult_vmat(3,0)(28)
		);


		FA_2_27_2: FA PORT MAP (
			mult_vmat(2,3)(27),
			mult_vmat(2,4)(27),
			mult_vmat(2,5)(27),
			mult_vmat(3,4)(27),
			mult_vmat(3,1)(28)
		);


		FA_2_27_3: FA PORT MAP (
			mult_vmat(2,6)(27),
			mult_vmat(2,7)(27),
			mult_vmat(2,8)(27),
			mult_vmat(3,5)(27),
			mult_vmat(3,2)(28)
		);


		-- COLUMN 29

		FA_2_28_1: FA PORT MAP (
			mult_vmat(2,0)(28),
			mult_vmat(2,1)(28),
			mult_vmat(2,2)(28),
			mult_vmat(3,3)(28),
			mult_vmat(3,0)(29)
		);


		FA_2_28_2: FA PORT MAP (
			mult_vmat(2,3)(28),
			mult_vmat(2,4)(28),
			mult_vmat(2,5)(28),
			mult_vmat(3,4)(28),
			mult_vmat(3,1)(29)
		);


		FA_2_28_3: FA PORT MAP (
			mult_vmat(2,6)(28),
			mult_vmat(2,7)(28),
			mult_vmat(2,8)(28),
			mult_vmat(3,5)(28),
			mult_vmat(3,2)(29)
		);


		-- COLUMN 30

		FA_2_29_1: FA PORT MAP (
			mult_vmat(2,0)(29),
			mult_vmat(2,1)(29),
			mult_vmat(2,2)(29),
			mult_vmat(3,3)(29),
			mult_vmat(3,0)(30)
		);


		FA_2_29_2: FA PORT MAP (
			mult_vmat(2,3)(29),
			mult_vmat(2,4)(29),
			mult_vmat(2,5)(29),
			mult_vmat(3,4)(29),
			mult_vmat(3,1)(30)
		);


		FA_2_29_3: FA PORT MAP (
			mult_vmat(2,6)(29),
			mult_vmat(2,7)(29),
			mult_vmat(2,8)(29),
			mult_vmat(3,5)(29),
			mult_vmat(3,2)(30)
		);


		-- COLUMN 31

		FA_2_30_1: FA PORT MAP (
			mult_vmat(2,0)(30),
			mult_vmat(2,1)(30),
			mult_vmat(2,2)(30),
			mult_vmat(3,3)(30),
			mult_vmat(3,0)(31)
		);


		FA_2_30_2: FA PORT MAP (
			mult_vmat(2,3)(30),
			mult_vmat(2,4)(30),
			mult_vmat(2,5)(30),
			mult_vmat(3,4)(30),
			mult_vmat(3,1)(31)
		);


		FA_2_30_3: FA PORT MAP (
			mult_vmat(2,6)(30),
			mult_vmat(2,7)(30),
			mult_vmat(2,8)(30),
			mult_vmat(3,5)(30),
			mult_vmat(3,2)(31)
		);


		-- COLUMN 32

		FA_2_31_1: FA PORT MAP (
			mult_vmat(2,0)(31),
			mult_vmat(2,1)(31),
			mult_vmat(2,2)(31),
			mult_vmat(3,3)(31),
			mult_vmat(3,0)(32)
		);


		FA_2_31_2: FA PORT MAP (
			mult_vmat(2,3)(31),
			mult_vmat(2,4)(31),
			mult_vmat(2,5)(31),
			mult_vmat(3,4)(31),
			mult_vmat(3,1)(32)
		);


		FA_2_31_3: FA PORT MAP (
			mult_vmat(2,6)(31),
			mult_vmat(2,7)(31),
			mult_vmat(2,8)(31),
			mult_vmat(3,5)(31),
			mult_vmat(3,2)(32)
		);


		-- COLUMN 33

		FA_2_32_1: FA PORT MAP (
			mult_vmat(2,0)(32),
			mult_vmat(2,1)(32),
			mult_vmat(2,2)(32),
			mult_vmat(3,3)(32),
			mult_vmat(3,0)(33)
		);


		FA_2_32_2: FA PORT MAP (
			mult_vmat(2,3)(32),
			mult_vmat(2,4)(32),
			mult_vmat(2,5)(32),
			mult_vmat(3,4)(32),
			mult_vmat(3,1)(33)
		);


		FA_2_32_3: FA PORT MAP (
			mult_vmat(2,6)(32),
			mult_vmat(2,7)(32),
			mult_vmat(2,8)(32),
			mult_vmat(3,5)(32),
			mult_vmat(3,2)(33)
		);


		-- COLUMN 34

		FA_2_33_1: FA PORT MAP (
			mult_vmat(2,0)(33),
			mult_vmat(2,1)(33),
			mult_vmat(2,2)(33),
			mult_vmat(3,3)(33),
			mult_vmat(3,0)(34)
		);


		FA_2_33_2: FA PORT MAP (
			mult_vmat(2,3)(33),
			mult_vmat(2,4)(33),
			mult_vmat(2,5)(33),
			mult_vmat(3,4)(33),
			mult_vmat(3,1)(34)
		);


		FA_2_33_3: FA PORT MAP (
			mult_vmat(2,6)(33),
			mult_vmat(2,7)(33),
			mult_vmat(2,8)(33),
			mult_vmat(3,5)(33),
			mult_vmat(3,2)(34)
		);


		-- COLUMN 35

		FA_2_34_1: FA PORT MAP (
			mult_vmat(2,0)(34),
			mult_vmat(2,1)(34),
			mult_vmat(2,2)(34),
			mult_vmat(3,3)(34),
			mult_vmat(3,0)(35)
		);


		FA_2_34_2: FA PORT MAP (
			mult_vmat(2,3)(34),
			mult_vmat(2,4)(34),
			mult_vmat(2,5)(34),
			mult_vmat(3,4)(34),
			mult_vmat(3,1)(35)
		);


		FA_2_34_3: FA PORT MAP (
			mult_vmat(2,6)(34),
			mult_vmat(2,7)(34),
			mult_vmat(2,8)(34),
			mult_vmat(3,5)(34),
			mult_vmat(3,2)(35)
		);


		-- COLUMN 36

		FA_2_35_1: FA PORT MAP (
			mult_vmat(2,0)(35),
			mult_vmat(2,1)(35),
			mult_vmat(2,2)(35),
			mult_vmat(3,3)(35),
			mult_vmat(3,0)(36)
		);


		FA_2_35_2: FA PORT MAP (
			mult_vmat(2,3)(35),
			mult_vmat(2,4)(35),
			mult_vmat(2,5)(35),
			mult_vmat(3,4)(35),
			mult_vmat(3,1)(36)
		);


		FA_2_35_3: FA PORT MAP (
			mult_vmat(2,6)(35),
			mult_vmat(2,7)(35),
			mult_vmat(2,8)(35),
			mult_vmat(3,5)(35),
			mult_vmat(3,2)(36)
		);


		-- COLUMN 37

		FA_2_36_1: FA PORT MAP (
			mult_vmat(2,0)(36),
			mult_vmat(2,1)(36),
			mult_vmat(2,2)(36),
			mult_vmat(3,3)(36),
			mult_vmat(3,0)(37)
		);


		FA_2_36_2: FA PORT MAP (
			mult_vmat(2,3)(36),
			mult_vmat(2,4)(36),
			mult_vmat(2,5)(36),
			mult_vmat(3,4)(36),
			mult_vmat(3,1)(37)
		);


		FA_2_36_3: FA PORT MAP (
			mult_vmat(2,6)(36),
			mult_vmat(2,7)(36),
			mult_vmat(2,8)(36),
			mult_vmat(3,5)(36),
			mult_vmat(3,2)(37)
		);


		-- COLUMN 38

		FA_2_37_1: FA PORT MAP (
			mult_vmat(2,0)(37),
			mult_vmat(2,1)(37),
			mult_vmat(2,2)(37),
			mult_vmat(3,3)(37),
			mult_vmat(3,0)(38)
		);


		FA_2_37_2: FA PORT MAP (
			mult_vmat(2,3)(37),
			mult_vmat(2,4)(37),
			mult_vmat(2,5)(37),
			mult_vmat(3,4)(37),
			mult_vmat(3,1)(38)
		);


		FA_2_37_3: FA PORT MAP (
			mult_vmat(2,6)(37),
			mult_vmat(2,7)(37),
			mult_vmat(2,8)(37),
			mult_vmat(3,5)(37),
			mult_vmat(3,2)(38)
		);


		-- COLUMN 39

		FA_2_38_1: FA PORT MAP (
			mult_vmat(2,0)(38),
			mult_vmat(2,1)(38),
			mult_vmat(2,2)(38),
			mult_vmat(3,3)(38),
			mult_vmat(3,0)(39)
		);


		FA_2_38_2: FA PORT MAP (
			mult_vmat(2,3)(38),
			mult_vmat(2,4)(38),
			mult_vmat(2,5)(38),
			mult_vmat(3,4)(38),
			mult_vmat(3,1)(39)
		);


		FA_2_38_3: FA PORT MAP (
			mult_vmat(2,6)(38),
			mult_vmat(2,7)(38),
			mult_vmat(2,8)(38),
			mult_vmat(3,5)(38),
			mult_vmat(3,2)(39)
		);


		-- COLUMN 40

		FA_2_39_1: FA PORT MAP (
			mult_vmat(2,0)(39),
			mult_vmat(2,1)(39),
			mult_vmat(2,2)(39),
			mult_vmat(3,3)(39),
			mult_vmat(3,0)(40)
		);


		FA_2_39_2: FA PORT MAP (
			mult_vmat(2,3)(39),
			mult_vmat(2,4)(39),
			mult_vmat(2,5)(39),
			mult_vmat(3,4)(39),
			mult_vmat(3,1)(40)
		);


		FA_2_39_3: FA PORT MAP (
			mult_vmat(2,6)(39),
			mult_vmat(2,7)(39),
			mult_vmat(2,8)(39),
			mult_vmat(3,5)(39),
			mult_vmat(3,2)(40)
		);


		-- COLUMN 41

		FA_2_40_1: FA PORT MAP (
			mult_vmat(2,0)(40),
			mult_vmat(2,1)(40),
			mult_vmat(2,2)(40),
			mult_vmat(3,3)(40),
			mult_vmat(3,0)(41)
		);


		FA_2_40_2: FA PORT MAP (
			mult_vmat(2,3)(40),
			mult_vmat(2,4)(40),
			mult_vmat(2,5)(40),
			mult_vmat(3,4)(40),
			mult_vmat(3,1)(41)
		);


		FA_2_40_3: FA PORT MAP (
			mult_vmat(2,6)(40),
			mult_vmat(2,7)(40),
			mult_vmat(2,8)(40),
			mult_vmat(3,5)(40),
			mult_vmat(3,2)(41)
		);


		-- COLUMN 42

		FA_2_41_1: FA PORT MAP (
			mult_vmat(2,0)(41),
			mult_vmat(2,1)(41),
			mult_vmat(2,2)(41),
			mult_vmat(3,3)(41),
			mult_vmat(3,0)(42)
		);


		FA_2_41_2: FA PORT MAP (
			mult_vmat(2,3)(41),
			mult_vmat(2,4)(41),
			mult_vmat(2,5)(41),
			mult_vmat(3,4)(41),
			mult_vmat(3,1)(42)
		);


		FA_2_41_3: FA PORT MAP (
			mult_vmat(2,6)(41),
			mult_vmat(2,7)(41),
			mult_vmat(2,8)(41),
			mult_vmat(3,5)(41),
			mult_vmat(3,2)(42)
		);


		-- COLUMN 43

		FA_2_42_1: FA PORT MAP (
			mult_vmat(2,0)(42),
			mult_vmat(2,1)(42),
			mult_vmat(2,2)(42),
			mult_vmat(3,3)(42),
			mult_vmat(3,0)(43)
		);


		FA_2_42_2: FA PORT MAP (
			mult_vmat(2,3)(42),
			mult_vmat(2,4)(42),
			mult_vmat(2,5)(42),
			mult_vmat(3,4)(42),
			mult_vmat(3,1)(43)
		);


		FA_2_42_3: FA PORT MAP (
			mult_vmat(2,6)(42),
			mult_vmat(2,7)(42),
			mult_vmat(2,8)(42),
			mult_vmat(3,5)(42),
			mult_vmat(3,2)(43)
		);


		-- COLUMN 44

		FA_2_43_1: FA PORT MAP (
			mult_vmat(2,0)(43),
			mult_vmat(2,1)(43),
			mult_vmat(2,2)(43),
			mult_vmat(3,3)(43),
			mult_vmat(3,0)(44)
		);


		FA_2_43_2: FA PORT MAP (
			mult_vmat(2,3)(43),
			mult_vmat(2,4)(43),
			mult_vmat(2,5)(43),
			mult_vmat(3,4)(43),
			mult_vmat(3,1)(44)
		);


		FA_2_43_3: FA PORT MAP (
			mult_vmat(2,6)(43),
			mult_vmat(2,7)(43),
			mult_vmat(2,8)(43),
			mult_vmat(3,5)(43),
			mult_vmat(3,2)(44)
		);


		-- COLUMN 45

		FA_2_44_1: FA PORT MAP (
			mult_vmat(2,0)(44),
			mult_vmat(2,1)(44),
			mult_vmat(2,2)(44),
			mult_vmat(3,3)(44),
			mult_vmat(3,0)(45)
		);


		FA_2_44_2: FA PORT MAP (
			mult_vmat(2,3)(44),
			mult_vmat(2,4)(44),
			mult_vmat(2,5)(44),
			mult_vmat(3,4)(44),
			mult_vmat(3,1)(45)
		);


		FA_2_44_3: FA PORT MAP (
			mult_vmat(2,6)(44),
			mult_vmat(2,7)(44),
			mult_vmat(2,8)(44),
			mult_vmat(3,5)(44),
			mult_vmat(3,2)(45)
		);


		-- COLUMN 46

		FA_2_45_1: FA PORT MAP (
			mult_vmat(2,0)(45),
			mult_vmat(2,1)(45),
			mult_vmat(2,2)(45),
			mult_vmat(3,3)(45),
			mult_vmat(3,0)(46)
		);


		FA_2_45_2: FA PORT MAP (
			mult_vmat(2,3)(45),
			mult_vmat(2,4)(45),
			mult_vmat(2,5)(45),
			mult_vmat(3,4)(45),
			mult_vmat(3,1)(46)
		);


		FA_2_45_3: FA PORT MAP (
			mult_vmat(2,6)(45),
			mult_vmat(2,7)(45),
			mult_vmat(2,8)(45),
			mult_vmat(3,5)(45),
			mult_vmat(3,2)(46)
		);


		-- COLUMN 47

		FA_2_46_1: FA PORT MAP (
			mult_vmat(2,0)(46),
			mult_vmat(2,1)(46),
			mult_vmat(2,2)(46),
			mult_vmat(3,3)(46),
			mult_vmat(3,0)(47)
		);


		FA_2_46_2: FA PORT MAP (
			mult_vmat(2,3)(46),
			mult_vmat(2,4)(46),
			mult_vmat(2,5)(46),
			mult_vmat(3,4)(46),
			mult_vmat(3,1)(47)
		);


		FA_2_46_3: FA PORT MAP (
			mult_vmat(2,6)(46),
			mult_vmat(2,7)(46),
			mult_vmat(2,8)(46),
			mult_vmat(3,5)(46),
			mult_vmat(3,2)(47)
		);


		-- COLUMN 48

		FA_2_47_1: FA PORT MAP (
			mult_vmat(2,0)(47),
			mult_vmat(2,1)(47),
			mult_vmat(2,2)(47),
			mult_vmat(3,3)(47),
			mult_vmat(3,0)(48)
		);


		FA_2_47_2: FA PORT MAP (
			mult_vmat(2,3)(47),
			mult_vmat(2,4)(47),
			mult_vmat(2,5)(47),
			mult_vmat(3,4)(47),
			mult_vmat(3,1)(48)
		);


		FA_2_47_3: FA PORT MAP (
			mult_vmat(2,6)(47),
			mult_vmat(2,7)(47),
			mult_vmat(2,8)(47),
			mult_vmat(3,5)(47),
			mult_vmat(3,2)(48)
		);


		-- COLUMN 49

		FA_2_48_1: FA PORT MAP (
			mult_vmat(2,0)(48),
			mult_vmat(2,1)(48),
			mult_vmat(2,2)(48),
			mult_vmat(3,3)(48),
			mult_vmat(3,0)(49)
		);


		FA_2_48_2: FA PORT MAP (
			mult_vmat(2,3)(48),
			mult_vmat(2,4)(48),
			mult_vmat(2,5)(48),
			mult_vmat(3,4)(48),
			mult_vmat(3,1)(49)
		);


		FA_2_48_3: FA PORT MAP (
			mult_vmat(2,6)(48),
			mult_vmat(2,7)(48),
			mult_vmat(2,8)(48),
			mult_vmat(3,5)(48),
			mult_vmat(3,2)(49)
		);


		-- COLUMN 50

		FA_2_49_1: FA PORT MAP (
			mult_vmat(2,0)(49),
			mult_vmat(2,1)(49),
			mult_vmat(2,2)(49),
			mult_vmat(3,3)(49),
			mult_vmat(3,0)(50)
		);


		FA_2_49_2: FA PORT MAP (
			mult_vmat(2,3)(49),
			mult_vmat(2,4)(49),
			mult_vmat(2,5)(49),
			mult_vmat(3,4)(49),
			mult_vmat(3,1)(50)
		);


		FA_2_49_3: FA PORT MAP (
			mult_vmat(2,6)(49),
			mult_vmat(2,7)(49),
			mult_vmat(2,8)(49),
			mult_vmat(3,5)(49),
			mult_vmat(3,2)(50)
		);


		-- COLUMN 51

		FA_2_50_1: FA PORT MAP (
			mult_vmat(2,0)(50),
			mult_vmat(2,1)(50),
			mult_vmat(2,2)(50),
			mult_vmat(3,3)(50),
			mult_vmat(3,0)(51)
		);


		FA_2_50_2: FA PORT MAP (
			mult_vmat(2,3)(50),
			mult_vmat(2,4)(50),
			mult_vmat(2,5)(50),
			mult_vmat(3,4)(50),
			mult_vmat(3,1)(51)
		);


		FA_2_50_3: FA PORT MAP (
			mult_vmat(2,6)(50),
			mult_vmat(2,7)(50),
			mult_vmat(2,8)(50),
			mult_vmat(3,5)(50),
			mult_vmat(3,2)(51)
		);


		-- COLUMN 52

		FA_2_51_1: FA PORT MAP (
			mult_vmat(2,0)(51),
			mult_vmat(2,1)(51),
			mult_vmat(2,2)(51),
			mult_vmat(3,3)(51),
			mult_vmat(3,0)(52)
		);


		FA_2_51_2: FA PORT MAP (
			mult_vmat(2,3)(51),
			mult_vmat(2,4)(51),
			mult_vmat(2,5)(51),
			mult_vmat(3,4)(51),
			mult_vmat(3,1)(52)
		);


		FA_2_51_3: FA PORT MAP (
			mult_vmat(2,6)(51),
			mult_vmat(2,7)(51),
			mult_vmat(2,8)(51),
			mult_vmat(3,5)(51),
			mult_vmat(3,2)(52)
		);


		-- COLUMN 53

		FA_2_52_1: FA PORT MAP (
			mult_vmat(2,0)(52),
			mult_vmat(2,1)(52),
			mult_vmat(2,2)(52),
			mult_vmat(3,3)(52),
			mult_vmat(3,0)(53)
		);


		FA_2_52_2: FA PORT MAP (
			mult_vmat(2,3)(52),
			mult_vmat(2,4)(52),
			mult_vmat(2,5)(52),
			mult_vmat(3,4)(52),
			mult_vmat(3,1)(53)
		);


		HA_2_52: HA PORT MAP (
			mult_vmat(2,6)(52),
			mult_vmat(2,7)(52),
			mult_vmat(3,5)(52),
			mult_vmat(3,2)(53)
		);


		-- COLUMN 54

		FA_2_53_1: FA PORT MAP (
			mult_vmat(2,0)(53),
			mult_vmat(2,1)(53),
			mult_vmat(2,2)(53),
			mult_vmat(3,3)(53),
			mult_vmat(3,0)(54)
		);


		FA_2_53_2: FA PORT MAP (
			mult_vmat(2,3)(53),
			mult_vmat(2,4)(53),
			mult_vmat(2,5)(53),
			mult_vmat(3,4)(53),
			mult_vmat(3,1)(54)
		);

		mult_vmat(3,5)(53) <= mult_vmat(2,6)(53);

		-- COLUMN 55

		FA_2_54_1: FA PORT MAP (
			mult_vmat(2,0)(54),
			mult_vmat(2,1)(54),
			mult_vmat(2,2)(54),
			mult_vmat(3,2)(54),
			mult_vmat(3,0)(55)
		);


		HA_2_54: HA PORT MAP (
			mult_vmat(2,3)(54),
			mult_vmat(2,4)(54),
			mult_vmat(3,3)(54),
			mult_vmat(3,1)(55)
		);

		mult_vmat(3,4)(54) <= mult_vmat(2,5)(54);
		mult_vmat(3,5)(54) <= mult_vmat(2,6)(54);

		-- COLUMN 56

		FA_2_55_1: FA PORT MAP (
			mult_vmat(2,0)(55),
			mult_vmat(2,1)(55),
			mult_vmat(2,2)(55),
			mult_vmat(3,2)(55),
			mult_vmat(3,0)(56)
		);

		mult_vmat(3,3)(55) <= mult_vmat(2,3)(55);
		mult_vmat(3,4)(55) <= mult_vmat(2,4)(55);
		mult_vmat(3,5)(55) <= mult_vmat(2,5)(55);

		-- COLUMN 57

		HA_2_56: HA PORT MAP (
			mult_vmat(2,0)(56),
			mult_vmat(2,1)(56),
			mult_vmat(3,1)(56),
			mult_vmat(3,0)(57)
		);

		mult_vmat(3,2)(56) <= mult_vmat(2,2)(56);
		mult_vmat(3,3)(56) <= mult_vmat(2,3)(56);
		mult_vmat(3,4)(56) <= mult_vmat(2,4)(56);
		mult_vmat(3,5)(56) <= mult_vmat(2,5)(56);

		-- COLUMN 58
		mult_vmat(3,1)(57) <= mult_vmat(2,0)(57);
		mult_vmat(3,2)(57) <= mult_vmat(2,1)(57);
		mult_vmat(3,3)(57) <= mult_vmat(2,2)(57);
		mult_vmat(3,4)(57) <= mult_vmat(2,3)(57);
		mult_vmat(3,5)(57) <= mult_vmat(2,4)(57);

		-- COLUMN 59
		mult_vmat(3,0)(58) <= mult_vmat(2,0)(58);
		mult_vmat(3,1)(58) <= mult_vmat(2,1)(58);
		mult_vmat(3,2)(58) <= mult_vmat(2,2)(58);
		mult_vmat(3,3)(58) <= mult_vmat(2,3)(58);
		mult_vmat(3,4)(58) <= mult_vmat(2,4)(58);

		-- COLUMN 60
		mult_vmat(3,0)(59) <= mult_vmat(2,0)(59);
		mult_vmat(3,1)(59) <= mult_vmat(2,1)(59);
		mult_vmat(3,2)(59) <= mult_vmat(2,2)(59);
		mult_vmat(3,3)(59) <= mult_vmat(2,3)(59);

		-- COLUMN 61
		mult_vmat(3,0)(60) <= mult_vmat(2,0)(60);
		mult_vmat(3,1)(60) <= mult_vmat(2,1)(60);
		mult_vmat(3,2)(60) <= mult_vmat(2,2)(60);
		mult_vmat(3,3)(60) <= mult_vmat(2,3)(60);

		-- COLUMN 62
		mult_vmat(3,0)(61) <= mult_vmat(2,0)(61);
		mult_vmat(3,1)(61) <= mult_vmat(2,1)(61);
		mult_vmat(3,2)(61) <= mult_vmat(2,2)(61);

		-- COLUMN 63
		mult_vmat(3,0)(62) <= mult_vmat(2,0)(62);
		mult_vmat(3,1)(62) <= mult_vmat(2,1)(62);
		mult_vmat(3,2)(62) <= mult_vmat(2,2)(62);

		-- COLUMN 64
		mult_vmat(3,0)(63) <= mult_vmat(2,0)(63);
		mult_vmat(3,1)(63) <= mult_vmat(2,1)(63);


	------------------------------------------
	-- LEVEL 4
	------------------------------------------


		-- COLUMN 1
		mult_vmat(4,0)(0) <= mult_vmat(3,0)(0);
		mult_vmat(4,1)(0) <= mult_vmat(3,1)(0);

		-- COLUMN 2
		mult_vmat(4,0)(1) <= mult_vmat(3,0)(1);

		-- COLUMN 3
		mult_vmat(4,0)(2) <= mult_vmat(3,0)(2);
		mult_vmat(4,1)(2) <= mult_vmat(3,1)(2);
		mult_vmat(4,2)(2) <= mult_vmat(3,2)(2);

		-- COLUMN 4
		mult_vmat(4,0)(3) <= mult_vmat(3,0)(3);
		mult_vmat(4,1)(3) <= mult_vmat(3,1)(3);

		-- COLUMN 5
		mult_vmat(4,0)(4) <= mult_vmat(3,0)(4);
		mult_vmat(4,1)(4) <= mult_vmat(3,1)(4);
		mult_vmat(4,2)(4) <= mult_vmat(3,2)(4);
		mult_vmat(4,3)(4) <= mult_vmat(3,3)(4);

		-- COLUMN 6
		mult_vmat(4,0)(5) <= mult_vmat(3,0)(5);
		mult_vmat(4,1)(5) <= mult_vmat(3,1)(5);
		mult_vmat(4,2)(5) <= mult_vmat(3,2)(5);

		-- COLUMN 7

		HA_3_6: HA PORT MAP (
			mult_vmat(3,0)(6),
			mult_vmat(3,1)(6),
			mult_vmat(4,0)(6),
			mult_vmat(4,0)(7)
		);

		mult_vmat(4,1)(6) <= mult_vmat(3,2)(6);
		mult_vmat(4,2)(6) <= mult_vmat(3,3)(6);
		mult_vmat(4,3)(6) <= mult_vmat(3,4)(6);

		-- COLUMN 8

		HA_3_7: HA PORT MAP (
			mult_vmat(3,0)(7),
			mult_vmat(3,1)(7),
			mult_vmat(4,1)(7),
			mult_vmat(4,0)(8)
		);

		mult_vmat(4,2)(7) <= mult_vmat(3,2)(7);
		mult_vmat(4,3)(7) <= mult_vmat(3,3)(7);

		-- COLUMN 9

		FA_3_8_1: FA PORT MAP (
			mult_vmat(3,0)(8),
			mult_vmat(3,1)(8),
			mult_vmat(3,2)(8),
			mult_vmat(4,1)(8),
			mult_vmat(4,0)(9)
		);


		HA_3_8: HA PORT MAP (
			mult_vmat(3,3)(8),
			mult_vmat(3,4)(8),
			mult_vmat(4,2)(8),
			mult_vmat(4,1)(9)
		);

		mult_vmat(4,3)(8) <= mult_vmat(3,5)(8);

		-- COLUMN 10

		FA_3_9_1: FA PORT MAP (
			mult_vmat(3,0)(9),
			mult_vmat(3,1)(9),
			mult_vmat(3,2)(9),
			mult_vmat(4,2)(9),
			mult_vmat(4,0)(10)
		);


		HA_3_9: HA PORT MAP (
			mult_vmat(3,3)(9),
			mult_vmat(3,4)(9),
			mult_vmat(4,3)(9),
			mult_vmat(4,1)(10)
		);


		-- COLUMN 11

		FA_3_10_1: FA PORT MAP (
			mult_vmat(3,0)(10),
			mult_vmat(3,1)(10),
			mult_vmat(3,2)(10),
			mult_vmat(4,2)(10),
			mult_vmat(4,0)(11)
		);


		FA_3_10_2: FA PORT MAP (
			mult_vmat(3,3)(10),
			mult_vmat(3,4)(10),
			mult_vmat(3,5)(10),
			mult_vmat(4,3)(10),
			mult_vmat(4,1)(11)
		);


		-- COLUMN 12

		FA_3_11_1: FA PORT MAP (
			mult_vmat(3,0)(11),
			mult_vmat(3,1)(11),
			mult_vmat(3,2)(11),
			mult_vmat(4,2)(11),
			mult_vmat(4,0)(12)
		);


		FA_3_11_2: FA PORT MAP (
			mult_vmat(3,3)(11),
			mult_vmat(3,4)(11),
			mult_vmat(3,5)(11),
			mult_vmat(4,3)(11),
			mult_vmat(4,1)(12)
		);


		-- COLUMN 13

		FA_3_12_1: FA PORT MAP (
			mult_vmat(3,0)(12),
			mult_vmat(3,1)(12),
			mult_vmat(3,2)(12),
			mult_vmat(4,2)(12),
			mult_vmat(4,0)(13)
		);


		FA_3_12_2: FA PORT MAP (
			mult_vmat(3,3)(12),
			mult_vmat(3,4)(12),
			mult_vmat(3,5)(12),
			mult_vmat(4,3)(12),
			mult_vmat(4,1)(13)
		);


		-- COLUMN 14

		FA_3_13_1: FA PORT MAP (
			mult_vmat(3,0)(13),
			mult_vmat(3,1)(13),
			mult_vmat(3,2)(13),
			mult_vmat(4,2)(13),
			mult_vmat(4,0)(14)
		);


		FA_3_13_2: FA PORT MAP (
			mult_vmat(3,3)(13),
			mult_vmat(3,4)(13),
			mult_vmat(3,5)(13),
			mult_vmat(4,3)(13),
			mult_vmat(4,1)(14)
		);


		-- COLUMN 15

		FA_3_14_1: FA PORT MAP (
			mult_vmat(3,0)(14),
			mult_vmat(3,1)(14),
			mult_vmat(3,2)(14),
			mult_vmat(4,2)(14),
			mult_vmat(4,0)(15)
		);


		FA_3_14_2: FA PORT MAP (
			mult_vmat(3,3)(14),
			mult_vmat(3,4)(14),
			mult_vmat(3,5)(14),
			mult_vmat(4,3)(14),
			mult_vmat(4,1)(15)
		);


		-- COLUMN 16

		FA_3_15_1: FA PORT MAP (
			mult_vmat(3,0)(15),
			mult_vmat(3,1)(15),
			mult_vmat(3,2)(15),
			mult_vmat(4,2)(15),
			mult_vmat(4,0)(16)
		);


		FA_3_15_2: FA PORT MAP (
			mult_vmat(3,3)(15),
			mult_vmat(3,4)(15),
			mult_vmat(3,5)(15),
			mult_vmat(4,3)(15),
			mult_vmat(4,1)(16)
		);


		-- COLUMN 17

		FA_3_16_1: FA PORT MAP (
			mult_vmat(3,0)(16),
			mult_vmat(3,1)(16),
			mult_vmat(3,2)(16),
			mult_vmat(4,2)(16),
			mult_vmat(4,0)(17)
		);


		FA_3_16_2: FA PORT MAP (
			mult_vmat(3,3)(16),
			mult_vmat(3,4)(16),
			mult_vmat(3,5)(16),
			mult_vmat(4,3)(16),
			mult_vmat(4,1)(17)
		);


		-- COLUMN 18

		FA_3_17_1: FA PORT MAP (
			mult_vmat(3,0)(17),
			mult_vmat(3,1)(17),
			mult_vmat(3,2)(17),
			mult_vmat(4,2)(17),
			mult_vmat(4,0)(18)
		);


		FA_3_17_2: FA PORT MAP (
			mult_vmat(3,3)(17),
			mult_vmat(3,4)(17),
			mult_vmat(3,5)(17),
			mult_vmat(4,3)(17),
			mult_vmat(4,1)(18)
		);


		-- COLUMN 19

		FA_3_18_1: FA PORT MAP (
			mult_vmat(3,0)(18),
			mult_vmat(3,1)(18),
			mult_vmat(3,2)(18),
			mult_vmat(4,2)(18),
			mult_vmat(4,0)(19)
		);


		FA_3_18_2: FA PORT MAP (
			mult_vmat(3,3)(18),
			mult_vmat(3,4)(18),
			mult_vmat(3,5)(18),
			mult_vmat(4,3)(18),
			mult_vmat(4,1)(19)
		);


		-- COLUMN 20

		FA_3_19_1: FA PORT MAP (
			mult_vmat(3,0)(19),
			mult_vmat(3,1)(19),
			mult_vmat(3,2)(19),
			mult_vmat(4,2)(19),
			mult_vmat(4,0)(20)
		);


		FA_3_19_2: FA PORT MAP (
			mult_vmat(3,3)(19),
			mult_vmat(3,4)(19),
			mult_vmat(3,5)(19),
			mult_vmat(4,3)(19),
			mult_vmat(4,1)(20)
		);


		-- COLUMN 21

		FA_3_20_1: FA PORT MAP (
			mult_vmat(3,0)(20),
			mult_vmat(3,1)(20),
			mult_vmat(3,2)(20),
			mult_vmat(4,2)(20),
			mult_vmat(4,0)(21)
		);


		FA_3_20_2: FA PORT MAP (
			mult_vmat(3,3)(20),
			mult_vmat(3,4)(20),
			mult_vmat(3,5)(20),
			mult_vmat(4,3)(20),
			mult_vmat(4,1)(21)
		);


		-- COLUMN 22

		FA_3_21_1: FA PORT MAP (
			mult_vmat(3,0)(21),
			mult_vmat(3,1)(21),
			mult_vmat(3,2)(21),
			mult_vmat(4,2)(21),
			mult_vmat(4,0)(22)
		);


		FA_3_21_2: FA PORT MAP (
			mult_vmat(3,3)(21),
			mult_vmat(3,4)(21),
			mult_vmat(3,5)(21),
			mult_vmat(4,3)(21),
			mult_vmat(4,1)(22)
		);


		-- COLUMN 23

		FA_3_22_1: FA PORT MAP (
			mult_vmat(3,0)(22),
			mult_vmat(3,1)(22),
			mult_vmat(3,2)(22),
			mult_vmat(4,2)(22),
			mult_vmat(4,0)(23)
		);


		FA_3_22_2: FA PORT MAP (
			mult_vmat(3,3)(22),
			mult_vmat(3,4)(22),
			mult_vmat(3,5)(22),
			mult_vmat(4,3)(22),
			mult_vmat(4,1)(23)
		);


		-- COLUMN 24

		FA_3_23_1: FA PORT MAP (
			mult_vmat(3,0)(23),
			mult_vmat(3,1)(23),
			mult_vmat(3,2)(23),
			mult_vmat(4,2)(23),
			mult_vmat(4,0)(24)
		);


		FA_3_23_2: FA PORT MAP (
			mult_vmat(3,3)(23),
			mult_vmat(3,4)(23),
			mult_vmat(3,5)(23),
			mult_vmat(4,3)(23),
			mult_vmat(4,1)(24)
		);


		-- COLUMN 25

		FA_3_24_1: FA PORT MAP (
			mult_vmat(3,0)(24),
			mult_vmat(3,1)(24),
			mult_vmat(3,2)(24),
			mult_vmat(4,2)(24),
			mult_vmat(4,0)(25)
		);


		FA_3_24_2: FA PORT MAP (
			mult_vmat(3,3)(24),
			mult_vmat(3,4)(24),
			mult_vmat(3,5)(24),
			mult_vmat(4,3)(24),
			mult_vmat(4,1)(25)
		);


		-- COLUMN 26

		FA_3_25_1: FA PORT MAP (
			mult_vmat(3,0)(25),
			mult_vmat(3,1)(25),
			mult_vmat(3,2)(25),
			mult_vmat(4,2)(25),
			mult_vmat(4,0)(26)
		);


		FA_3_25_2: FA PORT MAP (
			mult_vmat(3,3)(25),
			mult_vmat(3,4)(25),
			mult_vmat(3,5)(25),
			mult_vmat(4,3)(25),
			mult_vmat(4,1)(26)
		);


		-- COLUMN 27

		FA_3_26_1: FA PORT MAP (
			mult_vmat(3,0)(26),
			mult_vmat(3,1)(26),
			mult_vmat(3,2)(26),
			mult_vmat(4,2)(26),
			mult_vmat(4,0)(27)
		);


		FA_3_26_2: FA PORT MAP (
			mult_vmat(3,3)(26),
			mult_vmat(3,4)(26),
			mult_vmat(3,5)(26),
			mult_vmat(4,3)(26),
			mult_vmat(4,1)(27)
		);


		-- COLUMN 28

		FA_3_27_1: FA PORT MAP (
			mult_vmat(3,0)(27),
			mult_vmat(3,1)(27),
			mult_vmat(3,2)(27),
			mult_vmat(4,2)(27),
			mult_vmat(4,0)(28)
		);


		FA_3_27_2: FA PORT MAP (
			mult_vmat(3,3)(27),
			mult_vmat(3,4)(27),
			mult_vmat(3,5)(27),
			mult_vmat(4,3)(27),
			mult_vmat(4,1)(28)
		);


		-- COLUMN 29

		FA_3_28_1: FA PORT MAP (
			mult_vmat(3,0)(28),
			mult_vmat(3,1)(28),
			mult_vmat(3,2)(28),
			mult_vmat(4,2)(28),
			mult_vmat(4,0)(29)
		);


		FA_3_28_2: FA PORT MAP (
			mult_vmat(3,3)(28),
			mult_vmat(3,4)(28),
			mult_vmat(3,5)(28),
			mult_vmat(4,3)(28),
			mult_vmat(4,1)(29)
		);


		-- COLUMN 30

		FA_3_29_1: FA PORT MAP (
			mult_vmat(3,0)(29),
			mult_vmat(3,1)(29),
			mult_vmat(3,2)(29),
			mult_vmat(4,2)(29),
			mult_vmat(4,0)(30)
		);


		FA_3_29_2: FA PORT MAP (
			mult_vmat(3,3)(29),
			mult_vmat(3,4)(29),
			mult_vmat(3,5)(29),
			mult_vmat(4,3)(29),
			mult_vmat(4,1)(30)
		);


		-- COLUMN 31

		FA_3_30_1: FA PORT MAP (
			mult_vmat(3,0)(30),
			mult_vmat(3,1)(30),
			mult_vmat(3,2)(30),
			mult_vmat(4,2)(30),
			mult_vmat(4,0)(31)
		);


		FA_3_30_2: FA PORT MAP (
			mult_vmat(3,3)(30),
			mult_vmat(3,4)(30),
			mult_vmat(3,5)(30),
			mult_vmat(4,3)(30),
			mult_vmat(4,1)(31)
		);


		-- COLUMN 32

		FA_3_31_1: FA PORT MAP (
			mult_vmat(3,0)(31),
			mult_vmat(3,1)(31),
			mult_vmat(3,2)(31),
			mult_vmat(4,2)(31),
			mult_vmat(4,0)(32)
		);


		FA_3_31_2: FA PORT MAP (
			mult_vmat(3,3)(31),
			mult_vmat(3,4)(31),
			mult_vmat(3,5)(31),
			mult_vmat(4,3)(31),
			mult_vmat(4,1)(32)
		);


		-- COLUMN 33

		FA_3_32_1: FA PORT MAP (
			mult_vmat(3,0)(32),
			mult_vmat(3,1)(32),
			mult_vmat(3,2)(32),
			mult_vmat(4,2)(32),
			mult_vmat(4,0)(33)
		);


		FA_3_32_2: FA PORT MAP (
			mult_vmat(3,3)(32),
			mult_vmat(3,4)(32),
			mult_vmat(3,5)(32),
			mult_vmat(4,3)(32),
			mult_vmat(4,1)(33)
		);


		-- COLUMN 34

		FA_3_33_1: FA PORT MAP (
			mult_vmat(3,0)(33),
			mult_vmat(3,1)(33),
			mult_vmat(3,2)(33),
			mult_vmat(4,2)(33),
			mult_vmat(4,0)(34)
		);


		FA_3_33_2: FA PORT MAP (
			mult_vmat(3,3)(33),
			mult_vmat(3,4)(33),
			mult_vmat(3,5)(33),
			mult_vmat(4,3)(33),
			mult_vmat(4,1)(34)
		);


		-- COLUMN 35

		FA_3_34_1: FA PORT MAP (
			mult_vmat(3,0)(34),
			mult_vmat(3,1)(34),
			mult_vmat(3,2)(34),
			mult_vmat(4,2)(34),
			mult_vmat(4,0)(35)
		);


		FA_3_34_2: FA PORT MAP (
			mult_vmat(3,3)(34),
			mult_vmat(3,4)(34),
			mult_vmat(3,5)(34),
			mult_vmat(4,3)(34),
			mult_vmat(4,1)(35)
		);


		-- COLUMN 36

		FA_3_35_1: FA PORT MAP (
			mult_vmat(3,0)(35),
			mult_vmat(3,1)(35),
			mult_vmat(3,2)(35),
			mult_vmat(4,2)(35),
			mult_vmat(4,0)(36)
		);


		FA_3_35_2: FA PORT MAP (
			mult_vmat(3,3)(35),
			mult_vmat(3,4)(35),
			mult_vmat(3,5)(35),
			mult_vmat(4,3)(35),
			mult_vmat(4,1)(36)
		);


		-- COLUMN 37

		FA_3_36_1: FA PORT MAP (
			mult_vmat(3,0)(36),
			mult_vmat(3,1)(36),
			mult_vmat(3,2)(36),
			mult_vmat(4,2)(36),
			mult_vmat(4,0)(37)
		);


		FA_3_36_2: FA PORT MAP (
			mult_vmat(3,3)(36),
			mult_vmat(3,4)(36),
			mult_vmat(3,5)(36),
			mult_vmat(4,3)(36),
			mult_vmat(4,1)(37)
		);


		-- COLUMN 38

		FA_3_37_1: FA PORT MAP (
			mult_vmat(3,0)(37),
			mult_vmat(3,1)(37),
			mult_vmat(3,2)(37),
			mult_vmat(4,2)(37),
			mult_vmat(4,0)(38)
		);


		FA_3_37_2: FA PORT MAP (
			mult_vmat(3,3)(37),
			mult_vmat(3,4)(37),
			mult_vmat(3,5)(37),
			mult_vmat(4,3)(37),
			mult_vmat(4,1)(38)
		);


		-- COLUMN 39

		FA_3_38_1: FA PORT MAP (
			mult_vmat(3,0)(38),
			mult_vmat(3,1)(38),
			mult_vmat(3,2)(38),
			mult_vmat(4,2)(38),
			mult_vmat(4,0)(39)
		);


		FA_3_38_2: FA PORT MAP (
			mult_vmat(3,3)(38),
			mult_vmat(3,4)(38),
			mult_vmat(3,5)(38),
			mult_vmat(4,3)(38),
			mult_vmat(4,1)(39)
		);


		-- COLUMN 40

		FA_3_39_1: FA PORT MAP (
			mult_vmat(3,0)(39),
			mult_vmat(3,1)(39),
			mult_vmat(3,2)(39),
			mult_vmat(4,2)(39),
			mult_vmat(4,0)(40)
		);


		FA_3_39_2: FA PORT MAP (
			mult_vmat(3,3)(39),
			mult_vmat(3,4)(39),
			mult_vmat(3,5)(39),
			mult_vmat(4,3)(39),
			mult_vmat(4,1)(40)
		);


		-- COLUMN 41

		FA_3_40_1: FA PORT MAP (
			mult_vmat(3,0)(40),
			mult_vmat(3,1)(40),
			mult_vmat(3,2)(40),
			mult_vmat(4,2)(40),
			mult_vmat(4,0)(41)
		);


		FA_3_40_2: FA PORT MAP (
			mult_vmat(3,3)(40),
			mult_vmat(3,4)(40),
			mult_vmat(3,5)(40),
			mult_vmat(4,3)(40),
			mult_vmat(4,1)(41)
		);


		-- COLUMN 42

		FA_3_41_1: FA PORT MAP (
			mult_vmat(3,0)(41),
			mult_vmat(3,1)(41),
			mult_vmat(3,2)(41),
			mult_vmat(4,2)(41),
			mult_vmat(4,0)(42)
		);


		FA_3_41_2: FA PORT MAP (
			mult_vmat(3,3)(41),
			mult_vmat(3,4)(41),
			mult_vmat(3,5)(41),
			mult_vmat(4,3)(41),
			mult_vmat(4,1)(42)
		);


		-- COLUMN 43

		FA_3_42_1: FA PORT MAP (
			mult_vmat(3,0)(42),
			mult_vmat(3,1)(42),
			mult_vmat(3,2)(42),
			mult_vmat(4,2)(42),
			mult_vmat(4,0)(43)
		);


		FA_3_42_2: FA PORT MAP (
			mult_vmat(3,3)(42),
			mult_vmat(3,4)(42),
			mult_vmat(3,5)(42),
			mult_vmat(4,3)(42),
			mult_vmat(4,1)(43)
		);


		-- COLUMN 44

		FA_3_43_1: FA PORT MAP (
			mult_vmat(3,0)(43),
			mult_vmat(3,1)(43),
			mult_vmat(3,2)(43),
			mult_vmat(4,2)(43),
			mult_vmat(4,0)(44)
		);


		FA_3_43_2: FA PORT MAP (
			mult_vmat(3,3)(43),
			mult_vmat(3,4)(43),
			mult_vmat(3,5)(43),
			mult_vmat(4,3)(43),
			mult_vmat(4,1)(44)
		);


		-- COLUMN 45

		FA_3_44_1: FA PORT MAP (
			mult_vmat(3,0)(44),
			mult_vmat(3,1)(44),
			mult_vmat(3,2)(44),
			mult_vmat(4,2)(44),
			mult_vmat(4,0)(45)
		);


		FA_3_44_2: FA PORT MAP (
			mult_vmat(3,3)(44),
			mult_vmat(3,4)(44),
			mult_vmat(3,5)(44),
			mult_vmat(4,3)(44),
			mult_vmat(4,1)(45)
		);


		-- COLUMN 46

		FA_3_45_1: FA PORT MAP (
			mult_vmat(3,0)(45),
			mult_vmat(3,1)(45),
			mult_vmat(3,2)(45),
			mult_vmat(4,2)(45),
			mult_vmat(4,0)(46)
		);


		FA_3_45_2: FA PORT MAP (
			mult_vmat(3,3)(45),
			mult_vmat(3,4)(45),
			mult_vmat(3,5)(45),
			mult_vmat(4,3)(45),
			mult_vmat(4,1)(46)
		);


		-- COLUMN 47

		FA_3_46_1: FA PORT MAP (
			mult_vmat(3,0)(46),
			mult_vmat(3,1)(46),
			mult_vmat(3,2)(46),
			mult_vmat(4,2)(46),
			mult_vmat(4,0)(47)
		);


		FA_3_46_2: FA PORT MAP (
			mult_vmat(3,3)(46),
			mult_vmat(3,4)(46),
			mult_vmat(3,5)(46),
			mult_vmat(4,3)(46),
			mult_vmat(4,1)(47)
		);


		-- COLUMN 48

		FA_3_47_1: FA PORT MAP (
			mult_vmat(3,0)(47),
			mult_vmat(3,1)(47),
			mult_vmat(3,2)(47),
			mult_vmat(4,2)(47),
			mult_vmat(4,0)(48)
		);


		FA_3_47_2: FA PORT MAP (
			mult_vmat(3,3)(47),
			mult_vmat(3,4)(47),
			mult_vmat(3,5)(47),
			mult_vmat(4,3)(47),
			mult_vmat(4,1)(48)
		);


		-- COLUMN 49

		FA_3_48_1: FA PORT MAP (
			mult_vmat(3,0)(48),
			mult_vmat(3,1)(48),
			mult_vmat(3,2)(48),
			mult_vmat(4,2)(48),
			mult_vmat(4,0)(49)
		);


		FA_3_48_2: FA PORT MAP (
			mult_vmat(3,3)(48),
			mult_vmat(3,4)(48),
			mult_vmat(3,5)(48),
			mult_vmat(4,3)(48),
			mult_vmat(4,1)(49)
		);


		-- COLUMN 50

		FA_3_49_1: FA PORT MAP (
			mult_vmat(3,0)(49),
			mult_vmat(3,1)(49),
			mult_vmat(3,2)(49),
			mult_vmat(4,2)(49),
			mult_vmat(4,0)(50)
		);


		FA_3_49_2: FA PORT MAP (
			mult_vmat(3,3)(49),
			mult_vmat(3,4)(49),
			mult_vmat(3,5)(49),
			mult_vmat(4,3)(49),
			mult_vmat(4,1)(50)
		);


		-- COLUMN 51

		FA_3_50_1: FA PORT MAP (
			mult_vmat(3,0)(50),
			mult_vmat(3,1)(50),
			mult_vmat(3,2)(50),
			mult_vmat(4,2)(50),
			mult_vmat(4,0)(51)
		);


		FA_3_50_2: FA PORT MAP (
			mult_vmat(3,3)(50),
			mult_vmat(3,4)(50),
			mult_vmat(3,5)(50),
			mult_vmat(4,3)(50),
			mult_vmat(4,1)(51)
		);


		-- COLUMN 52

		FA_3_51_1: FA PORT MAP (
			mult_vmat(3,0)(51),
			mult_vmat(3,1)(51),
			mult_vmat(3,2)(51),
			mult_vmat(4,2)(51),
			mult_vmat(4,0)(52)
		);


		FA_3_51_2: FA PORT MAP (
			mult_vmat(3,3)(51),
			mult_vmat(3,4)(51),
			mult_vmat(3,5)(51),
			mult_vmat(4,3)(51),
			mult_vmat(4,1)(52)
		);


		-- COLUMN 53

		FA_3_52_1: FA PORT MAP (
			mult_vmat(3,0)(52),
			mult_vmat(3,1)(52),
			mult_vmat(3,2)(52),
			mult_vmat(4,2)(52),
			mult_vmat(4,0)(53)
		);


		FA_3_52_2: FA PORT MAP (
			mult_vmat(3,3)(52),
			mult_vmat(3,4)(52),
			mult_vmat(3,5)(52),
			mult_vmat(4,3)(52),
			mult_vmat(4,1)(53)
		);


		-- COLUMN 54

		FA_3_53_1: FA PORT MAP (
			mult_vmat(3,0)(53),
			mult_vmat(3,1)(53),
			mult_vmat(3,2)(53),
			mult_vmat(4,2)(53),
			mult_vmat(4,0)(54)
		);


		FA_3_53_2: FA PORT MAP (
			mult_vmat(3,3)(53),
			mult_vmat(3,4)(53),
			mult_vmat(3,5)(53),
			mult_vmat(4,3)(53),
			mult_vmat(4,1)(54)
		);


		-- COLUMN 55

		FA_3_54_1: FA PORT MAP (
			mult_vmat(3,0)(54),
			mult_vmat(3,1)(54),
			mult_vmat(3,2)(54),
			mult_vmat(4,2)(54),
			mult_vmat(4,0)(55)
		);


		FA_3_54_2: FA PORT MAP (
			mult_vmat(3,3)(54),
			mult_vmat(3,4)(54),
			mult_vmat(3,5)(54),
			mult_vmat(4,3)(54),
			mult_vmat(4,1)(55)
		);


		-- COLUMN 56

		FA_3_55_1: FA PORT MAP (
			mult_vmat(3,0)(55),
			mult_vmat(3,1)(55),
			mult_vmat(3,2)(55),
			mult_vmat(4,2)(55),
			mult_vmat(4,0)(56)
		);


		FA_3_55_2: FA PORT MAP (
			mult_vmat(3,3)(55),
			mult_vmat(3,4)(55),
			mult_vmat(3,5)(55),
			mult_vmat(4,3)(55),
			mult_vmat(4,1)(56)
		);


		-- COLUMN 57

		FA_3_56_1: FA PORT MAP (
			mult_vmat(3,0)(56),
			mult_vmat(3,1)(56),
			mult_vmat(3,2)(56),
			mult_vmat(4,2)(56),
			mult_vmat(4,0)(57)
		);


		FA_3_56_2: FA PORT MAP (
			mult_vmat(3,3)(56),
			mult_vmat(3,4)(56),
			mult_vmat(3,5)(56),
			mult_vmat(4,3)(56),
			mult_vmat(4,1)(57)
		);


		-- COLUMN 58

		FA_3_57_1: FA PORT MAP (
			mult_vmat(3,0)(57),
			mult_vmat(3,1)(57),
			mult_vmat(3,2)(57),
			mult_vmat(4,2)(57),
			mult_vmat(4,0)(58)
		);


		FA_3_57_2: FA PORT MAP (
			mult_vmat(3,3)(57),
			mult_vmat(3,4)(57),
			mult_vmat(3,5)(57),
			mult_vmat(4,3)(57),
			mult_vmat(4,1)(58)
		);


		-- COLUMN 59

		FA_3_58_1: FA PORT MAP (
			mult_vmat(3,0)(58),
			mult_vmat(3,1)(58),
			mult_vmat(3,2)(58),
			mult_vmat(4,2)(58),
			mult_vmat(4,0)(59)
		);


		HA_3_58: HA PORT MAP (
			mult_vmat(3,3)(58),
			mult_vmat(3,4)(58),
			mult_vmat(4,3)(58),
			mult_vmat(4,1)(59)
		);


		-- COLUMN 60

		FA_3_59_1: FA PORT MAP (
			mult_vmat(3,0)(59),
			mult_vmat(3,1)(59),
			mult_vmat(3,2)(59),
			mult_vmat(4,2)(59),
			mult_vmat(4,0)(60)
		);

		mult_vmat(4,3)(59) <= mult_vmat(3,3)(59);

		-- COLUMN 61

		HA_3_60: HA PORT MAP (
			mult_vmat(3,0)(60),
			mult_vmat(3,1)(60),
			mult_vmat(4,1)(60),
			mult_vmat(4,0)(61)
		);

		mult_vmat(4,2)(60) <= mult_vmat(3,2)(60);
		mult_vmat(4,3)(60) <= mult_vmat(3,3)(60);

		-- COLUMN 62
		mult_vmat(4,1)(61) <= mult_vmat(3,0)(61);
		mult_vmat(4,2)(61) <= mult_vmat(3,1)(61);
		mult_vmat(4,3)(61) <= mult_vmat(3,2)(61);

		-- COLUMN 63
		mult_vmat(4,0)(62) <= mult_vmat(3,0)(62);
		mult_vmat(4,1)(62) <= mult_vmat(3,1)(62);
		mult_vmat(4,2)(62) <= mult_vmat(3,2)(62);

		-- COLUMN 64
		mult_vmat(4,0)(63) <= mult_vmat(3,0)(63);
		mult_vmat(4,1)(63) <= mult_vmat(3,1)(63);


	------------------------------------------
	-- LEVEL 5
	------------------------------------------


		-- COLUMN 1
		mult_vmat(5,0)(0) <= mult_vmat(4,0)(0);
		mult_vmat(5,1)(0) <= mult_vmat(4,1)(0);

		-- COLUMN 2
		mult_vmat(5,0)(1) <= mult_vmat(4,0)(1);

		-- COLUMN 3
		mult_vmat(5,0)(2) <= mult_vmat(4,0)(2);
		mult_vmat(5,1)(2) <= mult_vmat(4,1)(2);
		mult_vmat(5,2)(2) <= mult_vmat(4,2)(2);

		-- COLUMN 4
		mult_vmat(5,0)(3) <= mult_vmat(4,0)(3);
		mult_vmat(5,1)(3) <= mult_vmat(4,1)(3);

		-- COLUMN 5

		HA_4_4: HA PORT MAP (
			mult_vmat(4,0)(4),
			mult_vmat(4,1)(4),
			mult_vmat(5,0)(4),
			mult_vmat(5,0)(5)
		);

		mult_vmat(5,1)(4) <= mult_vmat(4,2)(4);
		mult_vmat(5,2)(4) <= mult_vmat(4,3)(4);

		-- COLUMN 6

		HA_4_5: HA PORT MAP (
			mult_vmat(4,0)(5),
			mult_vmat(4,1)(5),
			mult_vmat(5,1)(5),
			mult_vmat(5,0)(6)
		);

		mult_vmat(5,2)(5) <= mult_vmat(4,2)(5);

		-- COLUMN 7

		FA_4_6_1: FA PORT MAP (
			mult_vmat(4,0)(6),
			mult_vmat(4,1)(6),
			mult_vmat(4,2)(6),
			mult_vmat(5,1)(6),
			mult_vmat(5,0)(7)
		);

		mult_vmat(5,2)(6) <= mult_vmat(4,3)(6);

		-- COLUMN 8

		FA_4_7_1: FA PORT MAP (
			mult_vmat(4,0)(7),
			mult_vmat(4,1)(7),
			mult_vmat(4,2)(7),
			mult_vmat(5,1)(7),
			mult_vmat(5,0)(8)
		);

		mult_vmat(5,2)(7) <= mult_vmat(4,3)(7);

		-- COLUMN 9

		FA_4_8_1: FA PORT MAP (
			mult_vmat(4,0)(8),
			mult_vmat(4,1)(8),
			mult_vmat(4,2)(8),
			mult_vmat(5,1)(8),
			mult_vmat(5,0)(9)
		);

		mult_vmat(5,2)(8) <= mult_vmat(4,3)(8);

		-- COLUMN 10

		FA_4_9_1: FA PORT MAP (
			mult_vmat(4,0)(9),
			mult_vmat(4,1)(9),
			mult_vmat(4,2)(9),
			mult_vmat(5,1)(9),
			mult_vmat(5,0)(10)
		);

		mult_vmat(5,2)(9) <= mult_vmat(4,3)(9);

		-- COLUMN 11

		FA_4_10_1: FA PORT MAP (
			mult_vmat(4,0)(10),
			mult_vmat(4,1)(10),
			mult_vmat(4,2)(10),
			mult_vmat(5,1)(10),
			mult_vmat(5,0)(11)
		);

		mult_vmat(5,2)(10) <= mult_vmat(4,3)(10);

		-- COLUMN 12

		FA_4_11_1: FA PORT MAP (
			mult_vmat(4,0)(11),
			mult_vmat(4,1)(11),
			mult_vmat(4,2)(11),
			mult_vmat(5,1)(11),
			mult_vmat(5,0)(12)
		);

		mult_vmat(5,2)(11) <= mult_vmat(4,3)(11);

		-- COLUMN 13

		FA_4_12_1: FA PORT MAP (
			mult_vmat(4,0)(12),
			mult_vmat(4,1)(12),
			mult_vmat(4,2)(12),
			mult_vmat(5,1)(12),
			mult_vmat(5,0)(13)
		);

		mult_vmat(5,2)(12) <= mult_vmat(4,3)(12);

		-- COLUMN 14

		FA_4_13_1: FA PORT MAP (
			mult_vmat(4,0)(13),
			mult_vmat(4,1)(13),
			mult_vmat(4,2)(13),
			mult_vmat(5,1)(13),
			mult_vmat(5,0)(14)
		);

		mult_vmat(5,2)(13) <= mult_vmat(4,3)(13);

		-- COLUMN 15

		FA_4_14_1: FA PORT MAP (
			mult_vmat(4,0)(14),
			mult_vmat(4,1)(14),
			mult_vmat(4,2)(14),
			mult_vmat(5,1)(14),
			mult_vmat(5,0)(15)
		);

		mult_vmat(5,2)(14) <= mult_vmat(4,3)(14);

		-- COLUMN 16

		FA_4_15_1: FA PORT MAP (
			mult_vmat(4,0)(15),
			mult_vmat(4,1)(15),
			mult_vmat(4,2)(15),
			mult_vmat(5,1)(15),
			mult_vmat(5,0)(16)
		);

		mult_vmat(5,2)(15) <= mult_vmat(4,3)(15);

		-- COLUMN 17

		FA_4_16_1: FA PORT MAP (
			mult_vmat(4,0)(16),
			mult_vmat(4,1)(16),
			mult_vmat(4,2)(16),
			mult_vmat(5,1)(16),
			mult_vmat(5,0)(17)
		);

		mult_vmat(5,2)(16) <= mult_vmat(4,3)(16);

		-- COLUMN 18

		FA_4_17_1: FA PORT MAP (
			mult_vmat(4,0)(17),
			mult_vmat(4,1)(17),
			mult_vmat(4,2)(17),
			mult_vmat(5,1)(17),
			mult_vmat(5,0)(18)
		);

		mult_vmat(5,2)(17) <= mult_vmat(4,3)(17);

		-- COLUMN 19

		FA_4_18_1: FA PORT MAP (
			mult_vmat(4,0)(18),
			mult_vmat(4,1)(18),
			mult_vmat(4,2)(18),
			mult_vmat(5,1)(18),
			mult_vmat(5,0)(19)
		);

		mult_vmat(5,2)(18) <= mult_vmat(4,3)(18);

		-- COLUMN 20

		FA_4_19_1: FA PORT MAP (
			mult_vmat(4,0)(19),
			mult_vmat(4,1)(19),
			mult_vmat(4,2)(19),
			mult_vmat(5,1)(19),
			mult_vmat(5,0)(20)
		);

		mult_vmat(5,2)(19) <= mult_vmat(4,3)(19);

		-- COLUMN 21

		FA_4_20_1: FA PORT MAP (
			mult_vmat(4,0)(20),
			mult_vmat(4,1)(20),
			mult_vmat(4,2)(20),
			mult_vmat(5,1)(20),
			mult_vmat(5,0)(21)
		);

		mult_vmat(5,2)(20) <= mult_vmat(4,3)(20);

		-- COLUMN 22

		FA_4_21_1: FA PORT MAP (
			mult_vmat(4,0)(21),
			mult_vmat(4,1)(21),
			mult_vmat(4,2)(21),
			mult_vmat(5,1)(21),
			mult_vmat(5,0)(22)
		);

		mult_vmat(5,2)(21) <= mult_vmat(4,3)(21);

		-- COLUMN 23

		FA_4_22_1: FA PORT MAP (
			mult_vmat(4,0)(22),
			mult_vmat(4,1)(22),
			mult_vmat(4,2)(22),
			mult_vmat(5,1)(22),
			mult_vmat(5,0)(23)
		);

		mult_vmat(5,2)(22) <= mult_vmat(4,3)(22);

		-- COLUMN 24

		FA_4_23_1: FA PORT MAP (
			mult_vmat(4,0)(23),
			mult_vmat(4,1)(23),
			mult_vmat(4,2)(23),
			mult_vmat(5,1)(23),
			mult_vmat(5,0)(24)
		);

		mult_vmat(5,2)(23) <= mult_vmat(4,3)(23);

		-- COLUMN 25

		FA_4_24_1: FA PORT MAP (
			mult_vmat(4,0)(24),
			mult_vmat(4,1)(24),
			mult_vmat(4,2)(24),
			mult_vmat(5,1)(24),
			mult_vmat(5,0)(25)
		);

		mult_vmat(5,2)(24) <= mult_vmat(4,3)(24);

		-- COLUMN 26

		FA_4_25_1: FA PORT MAP (
			mult_vmat(4,0)(25),
			mult_vmat(4,1)(25),
			mult_vmat(4,2)(25),
			mult_vmat(5,1)(25),
			mult_vmat(5,0)(26)
		);

		mult_vmat(5,2)(25) <= mult_vmat(4,3)(25);

		-- COLUMN 27

		FA_4_26_1: FA PORT MAP (
			mult_vmat(4,0)(26),
			mult_vmat(4,1)(26),
			mult_vmat(4,2)(26),
			mult_vmat(5,1)(26),
			mult_vmat(5,0)(27)
		);

		mult_vmat(5,2)(26) <= mult_vmat(4,3)(26);

		-- COLUMN 28

		FA_4_27_1: FA PORT MAP (
			mult_vmat(4,0)(27),
			mult_vmat(4,1)(27),
			mult_vmat(4,2)(27),
			mult_vmat(5,1)(27),
			mult_vmat(5,0)(28)
		);

		mult_vmat(5,2)(27) <= mult_vmat(4,3)(27);

		-- COLUMN 29

		FA_4_28_1: FA PORT MAP (
			mult_vmat(4,0)(28),
			mult_vmat(4,1)(28),
			mult_vmat(4,2)(28),
			mult_vmat(5,1)(28),
			mult_vmat(5,0)(29)
		);

		mult_vmat(5,2)(28) <= mult_vmat(4,3)(28);

		-- COLUMN 30

		FA_4_29_1: FA PORT MAP (
			mult_vmat(4,0)(29),
			mult_vmat(4,1)(29),
			mult_vmat(4,2)(29),
			mult_vmat(5,1)(29),
			mult_vmat(5,0)(30)
		);

		mult_vmat(5,2)(29) <= mult_vmat(4,3)(29);

		-- COLUMN 31

		FA_4_30_1: FA PORT MAP (
			mult_vmat(4,0)(30),
			mult_vmat(4,1)(30),
			mult_vmat(4,2)(30),
			mult_vmat(5,1)(30),
			mult_vmat(5,0)(31)
		);

		mult_vmat(5,2)(30) <= mult_vmat(4,3)(30);

		-- COLUMN 32

		FA_4_31_1: FA PORT MAP (
			mult_vmat(4,0)(31),
			mult_vmat(4,1)(31),
			mult_vmat(4,2)(31),
			mult_vmat(5,1)(31),
			mult_vmat(5,0)(32)
		);

		mult_vmat(5,2)(31) <= mult_vmat(4,3)(31);

		-- COLUMN 33

		FA_4_32_1: FA PORT MAP (
			mult_vmat(4,0)(32),
			mult_vmat(4,1)(32),
			mult_vmat(4,2)(32),
			mult_vmat(5,1)(32),
			mult_vmat(5,0)(33)
		);

		mult_vmat(5,2)(32) <= mult_vmat(4,3)(32);

		-- COLUMN 34

		FA_4_33_1: FA PORT MAP (
			mult_vmat(4,0)(33),
			mult_vmat(4,1)(33),
			mult_vmat(4,2)(33),
			mult_vmat(5,1)(33),
			mult_vmat(5,0)(34)
		);

		mult_vmat(5,2)(33) <= mult_vmat(4,3)(33);

		-- COLUMN 35

		FA_4_34_1: FA PORT MAP (
			mult_vmat(4,0)(34),
			mult_vmat(4,1)(34),
			mult_vmat(4,2)(34),
			mult_vmat(5,1)(34),
			mult_vmat(5,0)(35)
		);

		mult_vmat(5,2)(34) <= mult_vmat(4,3)(34);

		-- COLUMN 36

		FA_4_35_1: FA PORT MAP (
			mult_vmat(4,0)(35),
			mult_vmat(4,1)(35),
			mult_vmat(4,2)(35),
			mult_vmat(5,1)(35),
			mult_vmat(5,0)(36)
		);

		mult_vmat(5,2)(35) <= mult_vmat(4,3)(35);

		-- COLUMN 37

		FA_4_36_1: FA PORT MAP (
			mult_vmat(4,0)(36),
			mult_vmat(4,1)(36),
			mult_vmat(4,2)(36),
			mult_vmat(5,1)(36),
			mult_vmat(5,0)(37)
		);

		mult_vmat(5,2)(36) <= mult_vmat(4,3)(36);

		-- COLUMN 38

		FA_4_37_1: FA PORT MAP (
			mult_vmat(4,0)(37),
			mult_vmat(4,1)(37),
			mult_vmat(4,2)(37),
			mult_vmat(5,1)(37),
			mult_vmat(5,0)(38)
		);

		mult_vmat(5,2)(37) <= mult_vmat(4,3)(37);

		-- COLUMN 39

		FA_4_38_1: FA PORT MAP (
			mult_vmat(4,0)(38),
			mult_vmat(4,1)(38),
			mult_vmat(4,2)(38),
			mult_vmat(5,1)(38),
			mult_vmat(5,0)(39)
		);

		mult_vmat(5,2)(38) <= mult_vmat(4,3)(38);

		-- COLUMN 40

		FA_4_39_1: FA PORT MAP (
			mult_vmat(4,0)(39),
			mult_vmat(4,1)(39),
			mult_vmat(4,2)(39),
			mult_vmat(5,1)(39),
			mult_vmat(5,0)(40)
		);

		mult_vmat(5,2)(39) <= mult_vmat(4,3)(39);

		-- COLUMN 41

		FA_4_40_1: FA PORT MAP (
			mult_vmat(4,0)(40),
			mult_vmat(4,1)(40),
			mult_vmat(4,2)(40),
			mult_vmat(5,1)(40),
			mult_vmat(5,0)(41)
		);

		mult_vmat(5,2)(40) <= mult_vmat(4,3)(40);

		-- COLUMN 42

		FA_4_41_1: FA PORT MAP (
			mult_vmat(4,0)(41),
			mult_vmat(4,1)(41),
			mult_vmat(4,2)(41),
			mult_vmat(5,1)(41),
			mult_vmat(5,0)(42)
		);

		mult_vmat(5,2)(41) <= mult_vmat(4,3)(41);

		-- COLUMN 43

		FA_4_42_1: FA PORT MAP (
			mult_vmat(4,0)(42),
			mult_vmat(4,1)(42),
			mult_vmat(4,2)(42),
			mult_vmat(5,1)(42),
			mult_vmat(5,0)(43)
		);

		mult_vmat(5,2)(42) <= mult_vmat(4,3)(42);

		-- COLUMN 44

		FA_4_43_1: FA PORT MAP (
			mult_vmat(4,0)(43),
			mult_vmat(4,1)(43),
			mult_vmat(4,2)(43),
			mult_vmat(5,1)(43),
			mult_vmat(5,0)(44)
		);

		mult_vmat(5,2)(43) <= mult_vmat(4,3)(43);

		-- COLUMN 45

		FA_4_44_1: FA PORT MAP (
			mult_vmat(4,0)(44),
			mult_vmat(4,1)(44),
			mult_vmat(4,2)(44),
			mult_vmat(5,1)(44),
			mult_vmat(5,0)(45)
		);

		mult_vmat(5,2)(44) <= mult_vmat(4,3)(44);

		-- COLUMN 46

		FA_4_45_1: FA PORT MAP (
			mult_vmat(4,0)(45),
			mult_vmat(4,1)(45),
			mult_vmat(4,2)(45),
			mult_vmat(5,1)(45),
			mult_vmat(5,0)(46)
		);

		mult_vmat(5,2)(45) <= mult_vmat(4,3)(45);

		-- COLUMN 47

		FA_4_46_1: FA PORT MAP (
			mult_vmat(4,0)(46),
			mult_vmat(4,1)(46),
			mult_vmat(4,2)(46),
			mult_vmat(5,1)(46),
			mult_vmat(5,0)(47)
		);

		mult_vmat(5,2)(46) <= mult_vmat(4,3)(46);

		-- COLUMN 48

		FA_4_47_1: FA PORT MAP (
			mult_vmat(4,0)(47),
			mult_vmat(4,1)(47),
			mult_vmat(4,2)(47),
			mult_vmat(5,1)(47),
			mult_vmat(5,0)(48)
		);

		mult_vmat(5,2)(47) <= mult_vmat(4,3)(47);

		-- COLUMN 49

		FA_4_48_1: FA PORT MAP (
			mult_vmat(4,0)(48),
			mult_vmat(4,1)(48),
			mult_vmat(4,2)(48),
			mult_vmat(5,1)(48),
			mult_vmat(5,0)(49)
		);

		mult_vmat(5,2)(48) <= mult_vmat(4,3)(48);

		-- COLUMN 50

		FA_4_49_1: FA PORT MAP (
			mult_vmat(4,0)(49),
			mult_vmat(4,1)(49),
			mult_vmat(4,2)(49),
			mult_vmat(5,1)(49),
			mult_vmat(5,0)(50)
		);

		mult_vmat(5,2)(49) <= mult_vmat(4,3)(49);

		-- COLUMN 51

		FA_4_50_1: FA PORT MAP (
			mult_vmat(4,0)(50),
			mult_vmat(4,1)(50),
			mult_vmat(4,2)(50),
			mult_vmat(5,1)(50),
			mult_vmat(5,0)(51)
		);

		mult_vmat(5,2)(50) <= mult_vmat(4,3)(50);

		-- COLUMN 52

		FA_4_51_1: FA PORT MAP (
			mult_vmat(4,0)(51),
			mult_vmat(4,1)(51),
			mult_vmat(4,2)(51),
			mult_vmat(5,1)(51),
			mult_vmat(5,0)(52)
		);

		mult_vmat(5,2)(51) <= mult_vmat(4,3)(51);

		-- COLUMN 53

		FA_4_52_1: FA PORT MAP (
			mult_vmat(4,0)(52),
			mult_vmat(4,1)(52),
			mult_vmat(4,2)(52),
			mult_vmat(5,1)(52),
			mult_vmat(5,0)(53)
		);

		mult_vmat(5,2)(52) <= mult_vmat(4,3)(52);

		-- COLUMN 54

		FA_4_53_1: FA PORT MAP (
			mult_vmat(4,0)(53),
			mult_vmat(4,1)(53),
			mult_vmat(4,2)(53),
			mult_vmat(5,1)(53),
			mult_vmat(5,0)(54)
		);

		mult_vmat(5,2)(53) <= mult_vmat(4,3)(53);

		-- COLUMN 55

		FA_4_54_1: FA PORT MAP (
			mult_vmat(4,0)(54),
			mult_vmat(4,1)(54),
			mult_vmat(4,2)(54),
			mult_vmat(5,1)(54),
			mult_vmat(5,0)(55)
		);

		mult_vmat(5,2)(54) <= mult_vmat(4,3)(54);

		-- COLUMN 56

		FA_4_55_1: FA PORT MAP (
			mult_vmat(4,0)(55),
			mult_vmat(4,1)(55),
			mult_vmat(4,2)(55),
			mult_vmat(5,1)(55),
			mult_vmat(5,0)(56)
		);

		mult_vmat(5,2)(55) <= mult_vmat(4,3)(55);

		-- COLUMN 57

		FA_4_56_1: FA PORT MAP (
			mult_vmat(4,0)(56),
			mult_vmat(4,1)(56),
			mult_vmat(4,2)(56),
			mult_vmat(5,1)(56),
			mult_vmat(5,0)(57)
		);

		mult_vmat(5,2)(56) <= mult_vmat(4,3)(56);

		-- COLUMN 58

		FA_4_57_1: FA PORT MAP (
			mult_vmat(4,0)(57),
			mult_vmat(4,1)(57),
			mult_vmat(4,2)(57),
			mult_vmat(5,1)(57),
			mult_vmat(5,0)(58)
		);

		mult_vmat(5,2)(57) <= mult_vmat(4,3)(57);

		-- COLUMN 59

		FA_4_58_1: FA PORT MAP (
			mult_vmat(4,0)(58),
			mult_vmat(4,1)(58),
			mult_vmat(4,2)(58),
			mult_vmat(5,1)(58),
			mult_vmat(5,0)(59)
		);

		mult_vmat(5,2)(58) <= mult_vmat(4,3)(58);

		-- COLUMN 60

		FA_4_59_1: FA PORT MAP (
			mult_vmat(4,0)(59),
			mult_vmat(4,1)(59),
			mult_vmat(4,2)(59),
			mult_vmat(5,1)(59),
			mult_vmat(5,0)(60)
		);

		mult_vmat(5,2)(59) <= mult_vmat(4,3)(59);

		-- COLUMN 61

		FA_4_60_1: FA PORT MAP (
			mult_vmat(4,0)(60),
			mult_vmat(4,1)(60),
			mult_vmat(4,2)(60),
			mult_vmat(5,1)(60),
			mult_vmat(5,0)(61)
		);

		mult_vmat(5,2)(60) <= mult_vmat(4,3)(60);

		-- COLUMN 62

		FA_4_61_1: FA PORT MAP (
			mult_vmat(4,0)(61),
			mult_vmat(4,1)(61),
			mult_vmat(4,2)(61),
			mult_vmat(5,1)(61),
			mult_vmat(5,0)(62)
		);

		mult_vmat(5,2)(61) <= mult_vmat(4,3)(61);

		-- COLUMN 63

		HA_4_62: HA PORT MAP (
			mult_vmat(4,0)(62),
			mult_vmat(4,1)(62),
			mult_vmat(5,1)(62),
			mult_vmat(5,0)(63)
		);

		mult_vmat(5,2)(62) <= mult_vmat(4,2)(62);

		-- COLUMN 64
		mult_vmat(5,1)(63) <= mult_vmat(4,0)(63);
		mult_vmat(5,2)(63) <= mult_vmat(4,1)(63);


	------------------------------------------
	-- LEVEL 6
	------------------------------------------


		-- COLUMN 1
		mult_vmat(6,0)(0) <= mult_vmat(5,0)(0);
		mult_vmat(6,1)(0) <= mult_vmat(5,1)(0);

		-- COLUMN 2
		mult_vmat(6,0)(1) <= mult_vmat(5,0)(1);

		-- COLUMN 3

		HA_5_2: HA PORT MAP (
			mult_vmat(5,0)(2),
			mult_vmat(5,1)(2),
			mult_vmat(6,0)(2),
			mult_vmat(6,0)(3)
		);

		mult_vmat(6,1)(2) <= mult_vmat(5,2)(2);

		-- COLUMN 4

		HA_5_3: HA PORT MAP (
			mult_vmat(5,0)(3),
			mult_vmat(5,1)(3),
			mult_vmat(6,1)(3),
			mult_vmat(6,0)(4)
		);


		-- COLUMN 5

		FA_5_4_1: FA PORT MAP (
			mult_vmat(5,0)(4),
			mult_vmat(5,1)(4),
			mult_vmat(5,2)(4),
			mult_vmat(6,1)(4),
			mult_vmat(6,0)(5)
		);


		-- COLUMN 6

		FA_5_5_1: FA PORT MAP (
			mult_vmat(5,0)(5),
			mult_vmat(5,1)(5),
			mult_vmat(5,2)(5),
			mult_vmat(6,1)(5),
			mult_vmat(6,0)(6)
		);


		-- COLUMN 7

		FA_5_6_1: FA PORT MAP (
			mult_vmat(5,0)(6),
			mult_vmat(5,1)(6),
			mult_vmat(5,2)(6),
			mult_vmat(6,1)(6),
			mult_vmat(6,0)(7)
		);


		-- COLUMN 8

		FA_5_7_1: FA PORT MAP (
			mult_vmat(5,0)(7),
			mult_vmat(5,1)(7),
			mult_vmat(5,2)(7),
			mult_vmat(6,1)(7),
			mult_vmat(6,0)(8)
		);


		-- COLUMN 9

		FA_5_8_1: FA PORT MAP (
			mult_vmat(5,0)(8),
			mult_vmat(5,1)(8),
			mult_vmat(5,2)(8),
			mult_vmat(6,1)(8),
			mult_vmat(6,0)(9)
		);


		-- COLUMN 10

		FA_5_9_1: FA PORT MAP (
			mult_vmat(5,0)(9),
			mult_vmat(5,1)(9),
			mult_vmat(5,2)(9),
			mult_vmat(6,1)(9),
			mult_vmat(6,0)(10)
		);


		-- COLUMN 11

		FA_5_10_1: FA PORT MAP (
			mult_vmat(5,0)(10),
			mult_vmat(5,1)(10),
			mult_vmat(5,2)(10),
			mult_vmat(6,1)(10),
			mult_vmat(6,0)(11)
		);


		-- COLUMN 12

		FA_5_11_1: FA PORT MAP (
			mult_vmat(5,0)(11),
			mult_vmat(5,1)(11),
			mult_vmat(5,2)(11),
			mult_vmat(6,1)(11),
			mult_vmat(6,0)(12)
		);


		-- COLUMN 13

		FA_5_12_1: FA PORT MAP (
			mult_vmat(5,0)(12),
			mult_vmat(5,1)(12),
			mult_vmat(5,2)(12),
			mult_vmat(6,1)(12),
			mult_vmat(6,0)(13)
		);


		-- COLUMN 14

		FA_5_13_1: FA PORT MAP (
			mult_vmat(5,0)(13),
			mult_vmat(5,1)(13),
			mult_vmat(5,2)(13),
			mult_vmat(6,1)(13),
			mult_vmat(6,0)(14)
		);


		-- COLUMN 15

		FA_5_14_1: FA PORT MAP (
			mult_vmat(5,0)(14),
			mult_vmat(5,1)(14),
			mult_vmat(5,2)(14),
			mult_vmat(6,1)(14),
			mult_vmat(6,0)(15)
		);


		-- COLUMN 16

		FA_5_15_1: FA PORT MAP (
			mult_vmat(5,0)(15),
			mult_vmat(5,1)(15),
			mult_vmat(5,2)(15),
			mult_vmat(6,1)(15),
			mult_vmat(6,0)(16)
		);


		-- COLUMN 17

		FA_5_16_1: FA PORT MAP (
			mult_vmat(5,0)(16),
			mult_vmat(5,1)(16),
			mult_vmat(5,2)(16),
			mult_vmat(6,1)(16),
			mult_vmat(6,0)(17)
		);


		-- COLUMN 18

		FA_5_17_1: FA PORT MAP (
			mult_vmat(5,0)(17),
			mult_vmat(5,1)(17),
			mult_vmat(5,2)(17),
			mult_vmat(6,1)(17),
			mult_vmat(6,0)(18)
		);


		-- COLUMN 19

		FA_5_18_1: FA PORT MAP (
			mult_vmat(5,0)(18),
			mult_vmat(5,1)(18),
			mult_vmat(5,2)(18),
			mult_vmat(6,1)(18),
			mult_vmat(6,0)(19)
		);


		-- COLUMN 20

		FA_5_19_1: FA PORT MAP (
			mult_vmat(5,0)(19),
			mult_vmat(5,1)(19),
			mult_vmat(5,2)(19),
			mult_vmat(6,1)(19),
			mult_vmat(6,0)(20)
		);


		-- COLUMN 21

		FA_5_20_1: FA PORT MAP (
			mult_vmat(5,0)(20),
			mult_vmat(5,1)(20),
			mult_vmat(5,2)(20),
			mult_vmat(6,1)(20),
			mult_vmat(6,0)(21)
		);


		-- COLUMN 22

		FA_5_21_1: FA PORT MAP (
			mult_vmat(5,0)(21),
			mult_vmat(5,1)(21),
			mult_vmat(5,2)(21),
			mult_vmat(6,1)(21),
			mult_vmat(6,0)(22)
		);


		-- COLUMN 23

		FA_5_22_1: FA PORT MAP (
			mult_vmat(5,0)(22),
			mult_vmat(5,1)(22),
			mult_vmat(5,2)(22),
			mult_vmat(6,1)(22),
			mult_vmat(6,0)(23)
		);


		-- COLUMN 24

		FA_5_23_1: FA PORT MAP (
			mult_vmat(5,0)(23),
			mult_vmat(5,1)(23),
			mult_vmat(5,2)(23),
			mult_vmat(6,1)(23),
			mult_vmat(6,0)(24)
		);


		-- COLUMN 25

		FA_5_24_1: FA PORT MAP (
			mult_vmat(5,0)(24),
			mult_vmat(5,1)(24),
			mult_vmat(5,2)(24),
			mult_vmat(6,1)(24),
			mult_vmat(6,0)(25)
		);


		-- COLUMN 26

		FA_5_25_1: FA PORT MAP (
			mult_vmat(5,0)(25),
			mult_vmat(5,1)(25),
			mult_vmat(5,2)(25),
			mult_vmat(6,1)(25),
			mult_vmat(6,0)(26)
		);


		-- COLUMN 27

		FA_5_26_1: FA PORT MAP (
			mult_vmat(5,0)(26),
			mult_vmat(5,1)(26),
			mult_vmat(5,2)(26),
			mult_vmat(6,1)(26),
			mult_vmat(6,0)(27)
		);


		-- COLUMN 28

		FA_5_27_1: FA PORT MAP (
			mult_vmat(5,0)(27),
			mult_vmat(5,1)(27),
			mult_vmat(5,2)(27),
			mult_vmat(6,1)(27),
			mult_vmat(6,0)(28)
		);


		-- COLUMN 29

		FA_5_28_1: FA PORT MAP (
			mult_vmat(5,0)(28),
			mult_vmat(5,1)(28),
			mult_vmat(5,2)(28),
			mult_vmat(6,1)(28),
			mult_vmat(6,0)(29)
		);


		-- COLUMN 30

		FA_5_29_1: FA PORT MAP (
			mult_vmat(5,0)(29),
			mult_vmat(5,1)(29),
			mult_vmat(5,2)(29),
			mult_vmat(6,1)(29),
			mult_vmat(6,0)(30)
		);


		-- COLUMN 31

		FA_5_30_1: FA PORT MAP (
			mult_vmat(5,0)(30),
			mult_vmat(5,1)(30),
			mult_vmat(5,2)(30),
			mult_vmat(6,1)(30),
			mult_vmat(6,0)(31)
		);


		-- COLUMN 32

		FA_5_31_1: FA PORT MAP (
			mult_vmat(5,0)(31),
			mult_vmat(5,1)(31),
			mult_vmat(5,2)(31),
			mult_vmat(6,1)(31),
			mult_vmat(6,0)(32)
		);


		-- COLUMN 33

		FA_5_32_1: FA PORT MAP (
			mult_vmat(5,0)(32),
			mult_vmat(5,1)(32),
			mult_vmat(5,2)(32),
			mult_vmat(6,1)(32),
			mult_vmat(6,0)(33)
		);


		-- COLUMN 34

		FA_5_33_1: FA PORT MAP (
			mult_vmat(5,0)(33),
			mult_vmat(5,1)(33),
			mult_vmat(5,2)(33),
			mult_vmat(6,1)(33),
			mult_vmat(6,0)(34)
		);


		-- COLUMN 35

		FA_5_34_1: FA PORT MAP (
			mult_vmat(5,0)(34),
			mult_vmat(5,1)(34),
			mult_vmat(5,2)(34),
			mult_vmat(6,1)(34),
			mult_vmat(6,0)(35)
		);


		-- COLUMN 36

		FA_5_35_1: FA PORT MAP (
			mult_vmat(5,0)(35),
			mult_vmat(5,1)(35),
			mult_vmat(5,2)(35),
			mult_vmat(6,1)(35),
			mult_vmat(6,0)(36)
		);


		-- COLUMN 37

		FA_5_36_1: FA PORT MAP (
			mult_vmat(5,0)(36),
			mult_vmat(5,1)(36),
			mult_vmat(5,2)(36),
			mult_vmat(6,1)(36),
			mult_vmat(6,0)(37)
		);


		-- COLUMN 38

		FA_5_37_1: FA PORT MAP (
			mult_vmat(5,0)(37),
			mult_vmat(5,1)(37),
			mult_vmat(5,2)(37),
			mult_vmat(6,1)(37),
			mult_vmat(6,0)(38)
		);


		-- COLUMN 39

		FA_5_38_1: FA PORT MAP (
			mult_vmat(5,0)(38),
			mult_vmat(5,1)(38),
			mult_vmat(5,2)(38),
			mult_vmat(6,1)(38),
			mult_vmat(6,0)(39)
		);


		-- COLUMN 40

		FA_5_39_1: FA PORT MAP (
			mult_vmat(5,0)(39),
			mult_vmat(5,1)(39),
			mult_vmat(5,2)(39),
			mult_vmat(6,1)(39),
			mult_vmat(6,0)(40)
		);


		-- COLUMN 41

		FA_5_40_1: FA PORT MAP (
			mult_vmat(5,0)(40),
			mult_vmat(5,1)(40),
			mult_vmat(5,2)(40),
			mult_vmat(6,1)(40),
			mult_vmat(6,0)(41)
		);


		-- COLUMN 42

		FA_5_41_1: FA PORT MAP (
			mult_vmat(5,0)(41),
			mult_vmat(5,1)(41),
			mult_vmat(5,2)(41),
			mult_vmat(6,1)(41),
			mult_vmat(6,0)(42)
		);


		-- COLUMN 43

		FA_5_42_1: FA PORT MAP (
			mult_vmat(5,0)(42),
			mult_vmat(5,1)(42),
			mult_vmat(5,2)(42),
			mult_vmat(6,1)(42),
			mult_vmat(6,0)(43)
		);


		-- COLUMN 44

		FA_5_43_1: FA PORT MAP (
			mult_vmat(5,0)(43),
			mult_vmat(5,1)(43),
			mult_vmat(5,2)(43),
			mult_vmat(6,1)(43),
			mult_vmat(6,0)(44)
		);


		-- COLUMN 45

		FA_5_44_1: FA PORT MAP (
			mult_vmat(5,0)(44),
			mult_vmat(5,1)(44),
			mult_vmat(5,2)(44),
			mult_vmat(6,1)(44),
			mult_vmat(6,0)(45)
		);


		-- COLUMN 46

		FA_5_45_1: FA PORT MAP (
			mult_vmat(5,0)(45),
			mult_vmat(5,1)(45),
			mult_vmat(5,2)(45),
			mult_vmat(6,1)(45),
			mult_vmat(6,0)(46)
		);


		-- COLUMN 47

		FA_5_46_1: FA PORT MAP (
			mult_vmat(5,0)(46),
			mult_vmat(5,1)(46),
			mult_vmat(5,2)(46),
			mult_vmat(6,1)(46),
			mult_vmat(6,0)(47)
		);


		-- COLUMN 48

		FA_5_47_1: FA PORT MAP (
			mult_vmat(5,0)(47),
			mult_vmat(5,1)(47),
			mult_vmat(5,2)(47),
			mult_vmat(6,1)(47),
			mult_vmat(6,0)(48)
		);


		-- COLUMN 49

		FA_5_48_1: FA PORT MAP (
			mult_vmat(5,0)(48),
			mult_vmat(5,1)(48),
			mult_vmat(5,2)(48),
			mult_vmat(6,1)(48),
			mult_vmat(6,0)(49)
		);


		-- COLUMN 50

		FA_5_49_1: FA PORT MAP (
			mult_vmat(5,0)(49),
			mult_vmat(5,1)(49),
			mult_vmat(5,2)(49),
			mult_vmat(6,1)(49),
			mult_vmat(6,0)(50)
		);


		-- COLUMN 51

		FA_5_50_1: FA PORT MAP (
			mult_vmat(5,0)(50),
			mult_vmat(5,1)(50),
			mult_vmat(5,2)(50),
			mult_vmat(6,1)(50),
			mult_vmat(6,0)(51)
		);


		-- COLUMN 52

		FA_5_51_1: FA PORT MAP (
			mult_vmat(5,0)(51),
			mult_vmat(5,1)(51),
			mult_vmat(5,2)(51),
			mult_vmat(6,1)(51),
			mult_vmat(6,0)(52)
		);


		-- COLUMN 53

		FA_5_52_1: FA PORT MAP (
			mult_vmat(5,0)(52),
			mult_vmat(5,1)(52),
			mult_vmat(5,2)(52),
			mult_vmat(6,1)(52),
			mult_vmat(6,0)(53)
		);


		-- COLUMN 54

		FA_5_53_1: FA PORT MAP (
			mult_vmat(5,0)(53),
			mult_vmat(5,1)(53),
			mult_vmat(5,2)(53),
			mult_vmat(6,1)(53),
			mult_vmat(6,0)(54)
		);


		-- COLUMN 55

		FA_5_54_1: FA PORT MAP (
			mult_vmat(5,0)(54),
			mult_vmat(5,1)(54),
			mult_vmat(5,2)(54),
			mult_vmat(6,1)(54),
			mult_vmat(6,0)(55)
		);


		-- COLUMN 56

		FA_5_55_1: FA PORT MAP (
			mult_vmat(5,0)(55),
			mult_vmat(5,1)(55),
			mult_vmat(5,2)(55),
			mult_vmat(6,1)(55),
			mult_vmat(6,0)(56)
		);


		-- COLUMN 57

		FA_5_56_1: FA PORT MAP (
			mult_vmat(5,0)(56),
			mult_vmat(5,1)(56),
			mult_vmat(5,2)(56),
			mult_vmat(6,1)(56),
			mult_vmat(6,0)(57)
		);


		-- COLUMN 58

		FA_5_57_1: FA PORT MAP (
			mult_vmat(5,0)(57),
			mult_vmat(5,1)(57),
			mult_vmat(5,2)(57),
			mult_vmat(6,1)(57),
			mult_vmat(6,0)(58)
		);


		-- COLUMN 59

		FA_5_58_1: FA PORT MAP (
			mult_vmat(5,0)(58),
			mult_vmat(5,1)(58),
			mult_vmat(5,2)(58),
			mult_vmat(6,1)(58),
			mult_vmat(6,0)(59)
		);


		-- COLUMN 60

		FA_5_59_1: FA PORT MAP (
			mult_vmat(5,0)(59),
			mult_vmat(5,1)(59),
			mult_vmat(5,2)(59),
			mult_vmat(6,1)(59),
			mult_vmat(6,0)(60)
		);


		-- COLUMN 61

		FA_5_60_1: FA PORT MAP (
			mult_vmat(5,0)(60),
			mult_vmat(5,1)(60),
			mult_vmat(5,2)(60),
			mult_vmat(6,1)(60),
			mult_vmat(6,0)(61)
		);


		-- COLUMN 62

		FA_5_61_1: FA PORT MAP (
			mult_vmat(5,0)(61),
			mult_vmat(5,1)(61),
			mult_vmat(5,2)(61),
			mult_vmat(6,1)(61),
			mult_vmat(6,0)(62)
		);


		-- COLUMN 63

		FA_5_62_1: FA PORT MAP (
			mult_vmat(5,0)(62),
			mult_vmat(5,1)(62),
			mult_vmat(5,2)(62),
			mult_vmat(6,1)(62),
			mult_vmat(6,0)(63)
		);


		-- COLUMN 64

		FA_5_63_1: FA PORT MAP (
			mult_vmat(5,0)(63),
			mult_vmat(5,1)(63),
			mult_vmat(5,2)(63),
			mult_vmat(6,1)(63),

			open
		);




	------------------------------------------
	-- OUTPUTS
	------------------------------------------

		data_out1 <= mult_vmat(nl-1,0);
		data_out2 <= mult_vmat(nl-1,1);

END structure;