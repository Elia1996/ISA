library verilog;
use verilog.vl_types.all;
entity mul_pipe_tb is
end mul_pipe_tb;
