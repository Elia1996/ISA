library verilog;
use verilog.vl_types.all;
entity IIR_filter_optimized is
    port(
        DIN             : in     vl_logic_vector(11 downto 0);
        CLK             : in     vl_logic;
        RST_n           : in     vl_logic;
        VIN             : in     vl_logic;
        DOUT            : out    vl_logic_vector(11 downto 0);
        VOUT            : out    vl_logic
    );
end IIR_filter_optimized;
